//Secret key is'0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_c1908" written by ABC on Tue Nov  1 16:09:44 2022

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110,
    G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146,
    G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478,
    G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104,
    G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140,
    G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472,
    G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n526_,
    new_n528_, new_n529_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n536_, new_n537_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n548_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n123_));
  NAND2_X1  g001(.A1(new_n123_), .A2(KEYINPUT21), .ZN(new_n124_));
  INV_X1    g002(.A(G125), .ZN(new_n125_));
  NAND2_X1  g003(.A1(new_n125_), .A2(G140), .ZN(new_n126_));
  OAI21_X1  g004(.A(new_n124_), .B1(KEYINPUT21), .B2(new_n126_), .ZN(new_n127_));
  INV_X1    g005(.A(G146), .ZN(new_n128_));
  NAND2_X1  g006(.A1(new_n127_), .A2(new_n128_), .ZN(new_n129_));
  OAI211_X1 g007(.A(new_n124_), .B(G146), .C1(KEYINPUT21), .C2(new_n126_), .ZN(new_n130_));
  NAND2_X1  g008(.A1(new_n129_), .A2(new_n130_), .ZN(new_n131_));
  XNOR2_X1  g009(.A(G119), .B(G128), .ZN(new_n132_));
  INV_X1    g010(.A(G110), .ZN(new_n133_));
  XNOR2_X1  g011(.A(new_n132_), .B(new_n133_), .ZN(new_n134_));
  INV_X1    g012(.A(new_n134_), .ZN(new_n135_));
  NAND2_X1  g013(.A1(new_n131_), .A2(new_n135_), .ZN(new_n136_));
  INV_X1    g014(.A(G953), .ZN(new_n137_));
  NAND2_X1  g015(.A1(new_n137_), .A2(KEYINPUT10), .ZN(new_n138_));
  INV_X1    g016(.A(KEYINPUT10), .ZN(new_n139_));
  NAND2_X1  g017(.A1(new_n139_), .A2(G953), .ZN(new_n140_));
  AND2_X1   g018(.A1(new_n138_), .A2(new_n140_), .ZN(new_n141_));
  NAND3_X1  g019(.A1(new_n141_), .A2(G221), .A3(G234), .ZN(new_n142_));
  XNOR2_X1  g020(.A(new_n142_), .B(G137), .ZN(new_n143_));
  INV_X1    g021(.A(G140), .ZN(new_n144_));
  NOR3_X1   g022(.A1(new_n125_), .A2(new_n144_), .A3(KEYINPUT23), .ZN(new_n145_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n146_));
  AOI21_X1  g024(.A(new_n146_), .B1(G125), .B2(G140), .ZN(new_n147_));
  OAI22_X1  g025(.A1(new_n145_), .A2(new_n147_), .B1(G125), .B2(G140), .ZN(new_n148_));
  NAND2_X1  g026(.A1(new_n148_), .A2(new_n128_), .ZN(new_n149_));
  NAND3_X1  g027(.A1(new_n130_), .A2(new_n149_), .A3(new_n134_), .ZN(new_n150_));
  NAND3_X1  g028(.A1(new_n136_), .A2(new_n143_), .A3(new_n150_), .ZN(new_n151_));
  XOR2_X1   g029(.A(new_n142_), .B(G137), .Z(new_n152_));
  AOI21_X1  g030(.A(new_n134_), .B1(new_n129_), .B2(new_n130_), .ZN(new_n153_));
  AND3_X1   g031(.A1(new_n130_), .A2(new_n149_), .A3(new_n134_), .ZN(new_n154_));
  OAI21_X1  g032(.A(new_n152_), .B1(new_n153_), .B2(new_n154_), .ZN(new_n155_));
  AOI21_X1  g033(.A(G902), .B1(new_n151_), .B2(new_n155_), .ZN(new_n156_));
  INV_X1    g034(.A(G217), .ZN(new_n157_));
  INV_X1    g035(.A(G902), .ZN(new_n158_));
  AOI21_X1  g036(.A(new_n157_), .B1(G234), .B2(new_n158_), .ZN(new_n159_));
  INV_X1    g037(.A(new_n159_), .ZN(new_n160_));
  OR3_X1    g038(.A1(new_n156_), .A2(KEYINPUT26), .A3(new_n160_), .ZN(new_n161_));
  NAND2_X1  g039(.A1(new_n151_), .A2(new_n155_), .ZN(new_n162_));
  NAND3_X1  g040(.A1(new_n162_), .A2(new_n158_), .A3(new_n160_), .ZN(new_n163_));
  OAI21_X1  g041(.A(KEYINPUT26), .B1(new_n156_), .B2(new_n160_), .ZN(new_n164_));
  NAND3_X1  g042(.A1(new_n161_), .A2(new_n163_), .A3(new_n164_), .ZN(new_n165_));
  INV_X1    g043(.A(G472), .ZN(new_n166_));
  INV_X1    g044(.A(KEYINPUT27), .ZN(new_n167_));
  INV_X1    g045(.A(G237), .ZN(new_n168_));
  NAND4_X1  g046(.A1(new_n141_), .A2(new_n167_), .A3(G210), .A4(new_n168_), .ZN(new_n169_));
  NAND4_X1  g047(.A1(new_n138_), .A2(new_n140_), .A3(G210), .A4(new_n168_), .ZN(new_n170_));
  NAND2_X1  g048(.A1(new_n170_), .A2(KEYINPUT27), .ZN(new_n171_));
  NAND3_X1  g049(.A1(new_n169_), .A2(G101), .A3(new_n171_), .ZN(new_n172_));
  INV_X1    g050(.A(new_n172_), .ZN(new_n173_));
  AOI21_X1  g051(.A(G101), .B1(new_n169_), .B2(new_n171_), .ZN(new_n174_));
  OAI21_X1  g052(.A(KEYINPUT28), .B1(new_n173_), .B2(new_n174_), .ZN(new_n175_));
  NAND2_X1  g053(.A1(new_n169_), .A2(new_n171_), .ZN(new_n176_));
  INV_X1    g054(.A(G101), .ZN(new_n177_));
  NAND2_X1  g055(.A1(new_n176_), .A2(new_n177_), .ZN(new_n178_));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n179_));
  NAND3_X1  g057(.A1(new_n178_), .A2(new_n179_), .A3(new_n172_), .ZN(new_n180_));
  NAND2_X1  g058(.A1(new_n175_), .A2(new_n180_), .ZN(new_n181_));
  INV_X1    g059(.A(G128), .ZN(new_n182_));
  AND2_X1   g060(.A1(G143), .A2(G146), .ZN(new_n183_));
  NOR2_X1   g061(.A1(G143), .A2(G146), .ZN(new_n184_));
  OAI21_X1  g062(.A(new_n182_), .B1(new_n183_), .B2(new_n184_), .ZN(new_n185_));
  NAND2_X1  g063(.A1(new_n185_), .A2(KEYINPUT2), .ZN(new_n186_));
  INV_X1    g064(.A(G143), .ZN(new_n187_));
  NAND2_X1  g065(.A1(new_n187_), .A2(new_n128_), .ZN(new_n188_));
  NAND2_X1  g066(.A1(G143), .A2(G146), .ZN(new_n189_));
  NAND3_X1  g067(.A1(new_n188_), .A2(G128), .A3(new_n189_), .ZN(new_n190_));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n191_));
  NAND2_X1  g069(.A1(new_n190_), .A2(new_n191_), .ZN(new_n192_));
  NAND4_X1  g070(.A1(new_n188_), .A2(KEYINPUT3), .A3(G128), .A4(new_n189_), .ZN(new_n193_));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n194_));
  OAI211_X1 g072(.A(new_n194_), .B(new_n182_), .C1(new_n183_), .C2(new_n184_), .ZN(new_n195_));
  NAND4_X1  g073(.A1(new_n186_), .A2(new_n192_), .A3(new_n193_), .A4(new_n195_), .ZN(new_n196_));
  XNOR2_X1  g074(.A(G134), .B(G137), .ZN(new_n197_));
  INV_X1    g075(.A(G131), .ZN(new_n198_));
  XNOR2_X1  g076(.A(new_n197_), .B(new_n198_), .ZN(new_n199_));
  NAND2_X1  g077(.A1(new_n196_), .A2(new_n199_), .ZN(new_n200_));
  XNOR2_X1  g078(.A(G116), .B(G119), .ZN(new_n201_));
  INV_X1    g079(.A(G113), .ZN(new_n202_));
  NAND2_X1  g080(.A1(new_n201_), .A2(new_n202_), .ZN(new_n203_));
  INV_X1    g081(.A(new_n201_), .ZN(new_n204_));
  NAND2_X1  g082(.A1(new_n204_), .A2(G113), .ZN(new_n205_));
  XNOR2_X1  g083(.A(new_n197_), .B(G131), .ZN(new_n206_));
  AND2_X1   g084(.A1(new_n185_), .A2(new_n190_), .ZN(new_n207_));
  NAND2_X1  g085(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND4_X1  g086(.A1(new_n200_), .A2(new_n203_), .A3(new_n205_), .A4(new_n208_), .ZN(new_n209_));
  NAND2_X1  g087(.A1(new_n200_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g088(.A1(new_n205_), .A2(new_n203_), .ZN(new_n211_));
  NAND2_X1  g089(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  AND3_X1   g090(.A1(new_n181_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g091(.A(new_n181_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n214_));
  OAI211_X1 g092(.A(new_n166_), .B(new_n158_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g093(.A(new_n158_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g094(.A1(new_n216_), .A2(G472), .ZN(new_n217_));
  AOI21_X1  g095(.A(new_n165_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g096(.A(G214), .B1(G237), .B2(G902), .ZN(new_n219_));
  XNOR2_X1  g097(.A(new_n219_), .B(KEYINPUT0), .ZN(new_n220_));
  OAI21_X1  g098(.A(G210), .B1(G237), .B2(G902), .ZN(new_n221_));
  XNOR2_X1  g099(.A(new_n221_), .B(KEYINPUT9), .ZN(new_n222_));
  NAND2_X1  g100(.A1(new_n185_), .A2(new_n190_), .ZN(new_n223_));
  NAND2_X1  g101(.A1(new_n223_), .A2(new_n125_), .ZN(new_n224_));
  OAI21_X1  g102(.A(new_n224_), .B1(new_n196_), .B2(new_n125_), .ZN(new_n225_));
  NAND2_X1  g103(.A1(new_n137_), .A2(G224), .ZN(new_n226_));
  XOR2_X1   g104(.A(new_n226_), .B(KEYINPUT1), .Z(new_n227_));
  OR3_X1    g105(.A1(new_n225_), .A2(KEYINPUT6), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g106(.A(KEYINPUT5), .B1(new_n204_), .B2(G113), .ZN(new_n229_));
  INV_X1    g107(.A(new_n229_), .ZN(new_n230_));
  AND2_X1   g108(.A1(G104), .A2(G107), .ZN(new_n231_));
  NOR2_X1   g109(.A1(G104), .A2(G107), .ZN(new_n232_));
  OAI21_X1  g110(.A(new_n177_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g111(.A(G104), .ZN(new_n234_));
  INV_X1    g112(.A(G107), .ZN(new_n235_));
  NAND2_X1  g113(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g114(.A1(G104), .A2(G107), .ZN(new_n237_));
  NAND3_X1  g115(.A1(new_n236_), .A2(G101), .A3(new_n237_), .ZN(new_n238_));
  AND2_X1   g116(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g117(.A1(new_n204_), .A2(KEYINPUT5), .A3(G113), .ZN(new_n240_));
  NAND4_X1  g118(.A1(new_n230_), .A2(new_n203_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g119(.A(G110), .B(G122), .ZN(new_n242_));
  NAND2_X1  g120(.A1(new_n233_), .A2(new_n238_), .ZN(new_n243_));
  NAND2_X1  g121(.A1(new_n211_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g122(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g123(.A(new_n227_), .B1(new_n225_), .B2(KEYINPUT6), .ZN(new_n246_));
  NAND3_X1  g124(.A1(new_n228_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g125(.A1(new_n240_), .A2(new_n203_), .ZN(new_n248_));
  OAI21_X1  g126(.A(new_n243_), .B1(new_n248_), .B2(new_n229_), .ZN(new_n249_));
  NAND2_X1  g127(.A1(new_n249_), .A2(KEYINPUT7), .ZN(new_n250_));
  INV_X1    g128(.A(KEYINPUT7), .ZN(new_n251_));
  OAI211_X1 g129(.A(new_n251_), .B(new_n243_), .C1(new_n248_), .C2(new_n229_), .ZN(new_n252_));
  NAND3_X1  g130(.A1(new_n250_), .A2(new_n252_), .A3(new_n241_), .ZN(new_n253_));
  INV_X1    g131(.A(new_n242_), .ZN(new_n254_));
  NAND2_X1  g132(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g133(.A(KEYINPUT8), .ZN(new_n256_));
  NAND2_X1  g134(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g135(.A1(new_n253_), .A2(KEYINPUT8), .A3(new_n254_), .ZN(new_n258_));
  AOI21_X1  g136(.A(new_n247_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  AND3_X1   g137(.A1(new_n225_), .A2(KEYINPUT4), .A3(new_n227_), .ZN(new_n260_));
  AOI21_X1  g138(.A(KEYINPUT4), .B1(new_n225_), .B2(new_n227_), .ZN(new_n261_));
  OAI22_X1  g139(.A1(new_n260_), .A2(new_n261_), .B1(new_n227_), .B2(new_n225_), .ZN(new_n262_));
  NAND2_X1  g140(.A1(new_n241_), .A2(new_n244_), .ZN(new_n263_));
  NAND2_X1  g141(.A1(new_n263_), .A2(new_n254_), .ZN(new_n264_));
  NAND2_X1  g142(.A1(new_n264_), .A2(new_n245_), .ZN(new_n265_));
  NAND2_X1  g143(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g144(.A1(new_n266_), .A2(new_n158_), .ZN(new_n267_));
  OAI21_X1  g145(.A(new_n222_), .B1(new_n259_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g146(.A(new_n247_), .ZN(new_n269_));
  INV_X1    g147(.A(new_n258_), .ZN(new_n270_));
  AOI21_X1  g148(.A(KEYINPUT8), .B1(new_n253_), .B2(new_n254_), .ZN(new_n271_));
  OAI21_X1  g149(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g150(.A(G902), .B1(new_n262_), .B2(new_n265_), .ZN(new_n273_));
  INV_X1    g151(.A(new_n222_), .ZN(new_n274_));
  NAND3_X1  g152(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g153(.A(new_n220_), .B1(new_n268_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g154(.A1(G234), .A2(G237), .ZN(new_n277_));
  NAND3_X1  g155(.A1(new_n141_), .A2(G952), .A3(new_n277_), .ZN(new_n278_));
  NOR2_X1   g156(.A1(new_n158_), .A2(new_n137_), .ZN(new_n279_));
  INV_X1    g157(.A(G898), .ZN(new_n280_));
  NAND3_X1  g158(.A1(new_n279_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n281_));
  NAND2_X1  g159(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g160(.A(G113), .B(G122), .ZN(new_n283_));
  XNOR2_X1  g161(.A(new_n283_), .B(G104), .ZN(new_n284_));
  AND3_X1   g162(.A1(new_n168_), .A2(new_n137_), .A3(G214), .ZN(new_n285_));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n286_));
  NAND2_X1  g164(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g165(.A1(new_n168_), .A2(new_n137_), .A3(G214), .ZN(new_n288_));
  NAND2_X1  g166(.A1(new_n288_), .A2(KEYINPUT22), .ZN(new_n289_));
  AOI21_X1  g167(.A(G143), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g168(.A1(new_n138_), .A2(new_n140_), .A3(G214), .A4(new_n168_), .ZN(new_n291_));
  NOR2_X1   g169(.A1(new_n291_), .A2(new_n187_), .ZN(new_n292_));
  OR3_X1    g170(.A1(new_n290_), .A2(new_n292_), .A3(G131), .ZN(new_n293_));
  NOR2_X1   g171(.A1(new_n285_), .A2(G143), .ZN(new_n294_));
  OAI21_X1  g172(.A(G131), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g173(.A(new_n149_), .B1(new_n128_), .B2(new_n123_), .ZN(new_n296_));
  AND3_X1   g174(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g175(.A(new_n291_), .B(new_n187_), .ZN(new_n298_));
  NAND2_X1  g176(.A1(new_n298_), .A2(G131), .ZN(new_n299_));
  AOI21_X1  g177(.A(new_n131_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g178(.A(new_n284_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g179(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n302_));
  INV_X1    g180(.A(new_n284_), .ZN(new_n303_));
  NOR3_X1   g181(.A1(new_n290_), .A2(new_n292_), .A3(G131), .ZN(new_n304_));
  AOI21_X1  g182(.A(new_n304_), .B1(G131), .B2(new_n298_), .ZN(new_n305_));
  OAI211_X1 g183(.A(new_n302_), .B(new_n303_), .C1(new_n305_), .C2(new_n131_), .ZN(new_n306_));
  NAND2_X1  g184(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g185(.A1(new_n307_), .A2(new_n158_), .ZN(new_n308_));
  NAND2_X1  g186(.A1(new_n308_), .A2(G475), .ZN(new_n309_));
  INV_X1    g187(.A(G478), .ZN(new_n310_));
  INV_X1    g188(.A(G234), .ZN(new_n311_));
  NOR3_X1   g189(.A1(new_n157_), .A2(new_n311_), .A3(G953), .ZN(new_n312_));
  INV_X1    g190(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g191(.A(G116), .B(G122), .ZN(new_n314_));
  NAND2_X1  g192(.A1(new_n314_), .A2(new_n235_), .ZN(new_n315_));
  INV_X1    g193(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g194(.A1(new_n314_), .A2(new_n235_), .ZN(new_n317_));
  NAND2_X1  g195(.A1(new_n182_), .A2(G143), .ZN(new_n318_));
  NAND2_X1  g196(.A1(new_n187_), .A2(G128), .ZN(new_n319_));
  NAND2_X1  g197(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  OAI22_X1  g198(.A1(new_n316_), .A2(new_n317_), .B1(G134), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g199(.A(KEYINPUT17), .ZN(new_n322_));
  NAND2_X1  g200(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g201(.A1(new_n187_), .A2(KEYINPUT17), .A3(G128), .ZN(new_n324_));
  AOI22_X1  g202(.A1(new_n323_), .A2(new_n324_), .B1(new_n182_), .B2(G143), .ZN(new_n325_));
  INV_X1    g203(.A(KEYINPUT18), .ZN(new_n326_));
  INV_X1    g204(.A(G134), .ZN(new_n327_));
  OR3_X1    g205(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g206(.A(new_n326_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n329_));
  AOI21_X1  g207(.A(new_n321_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g208(.A1(new_n317_), .A2(KEYINPUT20), .ZN(new_n331_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n332_));
  OAI21_X1  g210(.A(new_n332_), .B1(new_n314_), .B2(new_n235_), .ZN(new_n333_));
  NAND3_X1  g211(.A1(new_n331_), .A2(new_n315_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g212(.A1(new_n320_), .A2(G134), .ZN(new_n335_));
  OR2_X1    g213(.A1(new_n335_), .A2(KEYINPUT19), .ZN(new_n336_));
  NOR2_X1   g214(.A1(new_n320_), .A2(G134), .ZN(new_n337_));
  AOI21_X1  g215(.A(new_n337_), .B1(KEYINPUT19), .B2(new_n335_), .ZN(new_n338_));
  AOI21_X1  g216(.A(new_n334_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g217(.A(new_n313_), .B1(new_n330_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g218(.A(new_n321_), .ZN(new_n341_));
  INV_X1    g219(.A(new_n329_), .ZN(new_n342_));
  NOR3_X1   g220(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n343_));
  OAI21_X1  g221(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g222(.A1(new_n338_), .A2(new_n336_), .ZN(new_n345_));
  AOI21_X1  g223(.A(new_n316_), .B1(KEYINPUT20), .B2(new_n317_), .ZN(new_n346_));
  NAND3_X1  g224(.A1(new_n345_), .A2(new_n333_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g225(.A1(new_n344_), .A2(new_n347_), .A3(new_n312_), .ZN(new_n348_));
  NAND2_X1  g226(.A1(new_n340_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g227(.A(new_n310_), .B1(new_n349_), .B2(new_n158_), .ZN(new_n350_));
  AOI211_X1 g228(.A(G478), .B(G902), .C1(new_n340_), .C2(new_n348_), .ZN(new_n351_));
  NOR2_X1   g229(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g230(.A1(G475), .A2(G902), .ZN(new_n353_));
  AND2_X1   g231(.A1(new_n187_), .A2(KEYINPUT24), .ZN(new_n354_));
  OR2_X1    g232(.A1(new_n291_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g233(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n187_), .ZN(new_n356_));
  AOI21_X1  g234(.A(new_n198_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g235(.A(new_n130_), .B(new_n149_), .C1(new_n304_), .C2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g236(.A(new_n303_), .B1(new_n358_), .B2(new_n302_), .ZN(new_n359_));
  INV_X1    g237(.A(KEYINPUT25), .ZN(new_n360_));
  AND2_X1   g238(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g239(.A(new_n306_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n362_));
  OAI21_X1  g240(.A(new_n353_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AND4_X1   g241(.A1(new_n282_), .A2(new_n309_), .A3(new_n352_), .A4(new_n363_), .ZN(new_n364_));
  AND2_X1   g242(.A1(new_n276_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g243(.A(KEYINPUT11), .ZN(new_n366_));
  NAND3_X1  g244(.A1(new_n207_), .A2(new_n239_), .A3(new_n366_), .ZN(new_n367_));
  NAND4_X1  g245(.A1(new_n190_), .A2(new_n185_), .A3(new_n233_), .A4(new_n238_), .ZN(new_n368_));
  NAND2_X1  g246(.A1(new_n368_), .A2(KEYINPUT11), .ZN(new_n369_));
  NAND2_X1  g247(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g248(.A1(new_n196_), .A2(new_n243_), .ZN(new_n371_));
  NAND3_X1  g249(.A1(new_n370_), .A2(new_n206_), .A3(new_n371_), .ZN(new_n372_));
  AOI22_X1  g250(.A1(new_n190_), .A2(new_n185_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n373_));
  INV_X1    g251(.A(KEYINPUT13), .ZN(new_n374_));
  OAI21_X1  g252(.A(new_n368_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g253(.A1(new_n223_), .A2(new_n243_), .ZN(new_n376_));
  NOR2_X1   g254(.A1(new_n376_), .A2(KEYINPUT13), .ZN(new_n377_));
  OAI211_X1 g255(.A(KEYINPUT14), .B(new_n199_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n378_));
  INV_X1    g256(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g257(.A1(new_n376_), .A2(KEYINPUT13), .ZN(new_n380_));
  NAND2_X1  g258(.A1(new_n373_), .A2(new_n374_), .ZN(new_n381_));
  NAND3_X1  g259(.A1(new_n380_), .A2(new_n381_), .A3(new_n368_), .ZN(new_n382_));
  AOI21_X1  g260(.A(KEYINPUT14), .B1(new_n382_), .B2(new_n199_), .ZN(new_n383_));
  OAI21_X1  g261(.A(new_n372_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g262(.A1(new_n141_), .A2(G227), .ZN(new_n385_));
  XNOR2_X1  g263(.A(G110), .B(G140), .ZN(new_n386_));
  XNOR2_X1  g264(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g265(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g266(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g267(.A(new_n206_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n390_));
  INV_X1    g268(.A(new_n390_), .ZN(new_n391_));
  AND4_X1   g269(.A1(KEYINPUT12), .A2(new_n370_), .A3(new_n206_), .A4(new_n371_), .ZN(new_n392_));
  AOI22_X1  g270(.A1(new_n367_), .A2(new_n369_), .B1(new_n196_), .B2(new_n243_), .ZN(new_n393_));
  AOI21_X1  g271(.A(KEYINPUT12), .B1(new_n393_), .B2(new_n206_), .ZN(new_n394_));
  OAI211_X1 g272(.A(new_n387_), .B(new_n391_), .C1(new_n392_), .C2(new_n394_), .ZN(new_n395_));
  AOI211_X1 g273(.A(KEYINPUT15), .B(G902), .C1(new_n389_), .C2(new_n395_), .ZN(new_n396_));
  INV_X1    g274(.A(KEYINPUT15), .ZN(new_n397_));
  AND3_X1   g275(.A1(new_n370_), .A2(new_n206_), .A3(new_n371_), .ZN(new_n398_));
  OAI21_X1  g276(.A(new_n199_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n399_));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n400_));
  NAND2_X1  g278(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g279(.A(new_n398_), .B1(new_n401_), .B2(new_n378_), .ZN(new_n402_));
  OAI21_X1  g280(.A(new_n395_), .B1(new_n387_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g281(.A(new_n397_), .B1(new_n403_), .B2(new_n158_), .ZN(new_n404_));
  OAI21_X1  g282(.A(G469), .B1(new_n396_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g283(.A1(new_n402_), .A2(new_n387_), .ZN(new_n406_));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n407_));
  NAND2_X1  g285(.A1(new_n372_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g286(.A1(new_n393_), .A2(KEYINPUT12), .A3(new_n206_), .ZN(new_n409_));
  AOI21_X1  g287(.A(new_n390_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g288(.A(new_n406_), .B1(new_n387_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g289(.A(G469), .ZN(new_n412_));
  NAND3_X1  g290(.A1(new_n411_), .A2(new_n412_), .A3(new_n158_), .ZN(new_n413_));
  NAND2_X1  g291(.A1(new_n405_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g292(.A(G221), .B1(new_n311_), .B2(G902), .ZN(new_n415_));
  AOI21_X1  g293(.A(KEYINPUT16), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n417_));
  INV_X1    g295(.A(new_n415_), .ZN(new_n418_));
  AOI211_X1 g296(.A(new_n417_), .B(new_n418_), .C1(new_n405_), .C2(new_n413_), .ZN(new_n419_));
  OAI211_X1 g297(.A(new_n218_), .B(new_n365_), .C1(new_n416_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g298(.A1(new_n420_), .A2(KEYINPUT29), .ZN(new_n421_));
  NOR2_X1   g299(.A1(new_n402_), .A2(new_n387_), .ZN(new_n422_));
  AOI211_X1 g300(.A(new_n388_), .B(new_n390_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n423_));
  OAI21_X1  g301(.A(new_n158_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g302(.A1(new_n424_), .A2(KEYINPUT15), .ZN(new_n425_));
  NAND3_X1  g303(.A1(new_n403_), .A2(new_n397_), .A3(new_n158_), .ZN(new_n426_));
  AOI21_X1  g304(.A(new_n412_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g305(.A(new_n413_), .ZN(new_n428_));
  OAI21_X1  g306(.A(new_n415_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g307(.A1(new_n429_), .A2(new_n417_), .ZN(new_n430_));
  NAND3_X1  g308(.A1(new_n414_), .A2(KEYINPUT16), .A3(new_n415_), .ZN(new_n431_));
  NAND2_X1  g309(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n433_));
  NAND4_X1  g311(.A1(new_n432_), .A2(new_n433_), .A3(new_n218_), .A4(new_n365_), .ZN(new_n434_));
  NAND2_X1  g312(.A1(new_n421_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g313(.A(new_n435_), .B(G101), .ZN(G3));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n437_));
  NAND2_X1  g315(.A1(new_n351_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g316(.A1(new_n349_), .A2(new_n310_), .A3(new_n158_), .ZN(new_n439_));
  NAND2_X1  g317(.A1(new_n439_), .A2(KEYINPUT30), .ZN(new_n440_));
  AOI21_X1  g318(.A(new_n350_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g319(.A1(new_n309_), .A2(new_n363_), .ZN(new_n442_));
  NAND2_X1  g320(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g321(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g322(.A1(new_n444_), .A2(new_n282_), .ZN(new_n445_));
  NAND2_X1  g323(.A1(new_n217_), .A2(new_n215_), .ZN(new_n446_));
  NOR2_X1   g324(.A1(new_n446_), .A2(new_n165_), .ZN(new_n447_));
  NAND2_X1  g325(.A1(new_n447_), .A2(new_n276_), .ZN(new_n448_));
  AOI211_X1 g326(.A(new_n445_), .B(new_n448_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n449_));
  XNOR2_X1  g327(.A(new_n449_), .B(new_n234_), .ZN(G6));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n451_));
  AOI21_X1  g329(.A(new_n451_), .B1(new_n307_), .B2(new_n158_), .ZN(new_n452_));
  AOI211_X1 g330(.A(KEYINPUT31), .B(G902), .C1(new_n301_), .C2(new_n306_), .ZN(new_n453_));
  OAI21_X1  g331(.A(G475), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g332(.A(new_n352_), .ZN(new_n455_));
  NAND3_X1  g333(.A1(new_n454_), .A2(new_n363_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g334(.A(new_n282_), .ZN(new_n457_));
  NOR2_X1   g335(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g336(.A(new_n458_), .ZN(new_n459_));
  AOI211_X1 g337(.A(new_n448_), .B(new_n459_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n460_));
  XNOR2_X1  g338(.A(new_n460_), .B(G107), .ZN(new_n461_));
  XNOR2_X1  g339(.A(new_n461_), .B(KEYINPUT32), .ZN(G9));
  INV_X1    g340(.A(KEYINPUT34), .ZN(new_n463_));
  AOI21_X1  g341(.A(KEYINPUT33), .B1(new_n162_), .B2(new_n160_), .ZN(new_n464_));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n465_));
  AOI211_X1 g343(.A(new_n465_), .B(new_n159_), .C1(new_n151_), .C2(new_n155_), .ZN(new_n466_));
  OAI21_X1  g344(.A(new_n158_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  OR2_X1    g345(.A1(new_n156_), .A2(new_n160_), .ZN(new_n468_));
  NAND2_X1  g346(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g347(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g348(.A(new_n463_), .B1(new_n470_), .B2(new_n446_), .ZN(new_n471_));
  NAND4_X1  g349(.A1(new_n469_), .A2(KEYINPUT34), .A3(new_n217_), .A4(new_n215_), .ZN(new_n472_));
  NAND2_X1  g350(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g351(.A(new_n365_), .B(new_n473_), .C1(new_n416_), .C2(new_n419_), .ZN(new_n474_));
  NAND2_X1  g352(.A1(new_n474_), .A2(KEYINPUT35), .ZN(new_n475_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n476_));
  NAND4_X1  g354(.A1(new_n432_), .A2(new_n476_), .A3(new_n365_), .A4(new_n473_), .ZN(new_n477_));
  NAND2_X1  g355(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g356(.A(new_n478_), .B(G110), .ZN(G12));
  AOI22_X1  g357(.A1(new_n217_), .A2(new_n215_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n480_));
  INV_X1    g358(.A(G900), .ZN(new_n481_));
  NAND3_X1  g359(.A1(new_n279_), .A2(new_n481_), .A3(new_n277_), .ZN(new_n482_));
  AND2_X1   g360(.A1(new_n278_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g361(.A1(new_n456_), .A2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g362(.A1(new_n432_), .A2(new_n276_), .A3(new_n480_), .A4(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g363(.A(new_n485_), .B(G128), .ZN(G30));
  NAND2_X1  g364(.A1(new_n268_), .A2(new_n275_), .ZN(new_n487_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n488_));
  XNOR2_X1  g366(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  AOI21_X1  g367(.A(new_n352_), .B1(new_n309_), .B2(new_n363_), .ZN(new_n490_));
  INV_X1    g368(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g369(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g370(.A(new_n209_), .B(KEYINPUT37), .ZN(new_n493_));
  NAND2_X1  g371(.A1(new_n493_), .A2(new_n212_), .ZN(new_n494_));
  INV_X1    g372(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g373(.A(new_n214_), .B1(new_n495_), .B2(new_n181_), .ZN(new_n496_));
  NOR2_X1   g374(.A1(new_n496_), .A2(G902), .ZN(new_n497_));
  OAI21_X1  g375(.A(new_n215_), .B1(new_n497_), .B2(new_n166_), .ZN(new_n498_));
  INV_X1    g376(.A(new_n220_), .ZN(new_n499_));
  NAND2_X1  g377(.A1(new_n499_), .A2(new_n415_), .ZN(new_n500_));
  NOR2_X1   g378(.A1(new_n483_), .A2(new_n500_), .ZN(new_n501_));
  AND4_X1   g379(.A1(new_n414_), .A2(new_n498_), .A3(new_n470_), .A4(new_n501_), .ZN(new_n502_));
  NAND2_X1  g380(.A1(new_n492_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g381(.A(new_n503_), .B(KEYINPUT38), .ZN(new_n504_));
  XNOR2_X1  g382(.A(new_n504_), .B(new_n187_), .ZN(G45));
  NOR2_X1   g383(.A1(new_n443_), .A2(new_n483_), .ZN(new_n506_));
  INV_X1    g384(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g385(.A1(new_n259_), .A2(new_n267_), .A3(new_n222_), .ZN(new_n508_));
  AOI21_X1  g386(.A(new_n274_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n509_));
  OAI21_X1  g387(.A(new_n499_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g388(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g389(.A1(new_n432_), .A2(new_n480_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g390(.A(new_n512_), .B(G146), .ZN(G48));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n514_));
  NAND2_X1  g392(.A1(new_n413_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g393(.A1(new_n411_), .A2(new_n158_), .ZN(new_n516_));
  NAND2_X1  g394(.A1(new_n516_), .A2(G469), .ZN(new_n517_));
  NAND4_X1  g395(.A1(new_n411_), .A2(KEYINPUT39), .A3(new_n412_), .A4(new_n158_), .ZN(new_n518_));
  NAND4_X1  g396(.A1(new_n515_), .A2(new_n517_), .A3(new_n415_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g397(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g398(.A(new_n165_), .ZN(new_n521_));
  NAND2_X1  g399(.A1(new_n521_), .A2(new_n446_), .ZN(new_n522_));
  NOR2_X1   g400(.A1(new_n510_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g401(.A1(new_n520_), .A2(new_n523_), .A3(new_n282_), .A4(new_n444_), .ZN(new_n524_));
  XNOR2_X1  g402(.A(new_n524_), .B(G113), .ZN(G15));
  NAND3_X1  g403(.A1(new_n520_), .A2(new_n523_), .A3(new_n458_), .ZN(new_n526_));
  XNOR2_X1  g404(.A(new_n526_), .B(G116), .ZN(G18));
  AND3_X1   g405(.A1(new_n276_), .A2(new_n364_), .A3(new_n480_), .ZN(new_n528_));
  NAND2_X1  g406(.A1(new_n528_), .A2(new_n520_), .ZN(new_n529_));
  XNOR2_X1  g407(.A(new_n529_), .B(G119), .ZN(G21));
  AND3_X1   g408(.A1(new_n515_), .A2(new_n518_), .A3(new_n517_), .ZN(new_n531_));
  AND2_X1   g409(.A1(new_n487_), .A2(new_n490_), .ZN(new_n532_));
  NOR4_X1   g410(.A1(new_n446_), .A2(new_n165_), .A3(new_n220_), .A4(new_n457_), .ZN(new_n533_));
  NAND4_X1  g411(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .A4(new_n415_), .ZN(new_n534_));
  XNOR2_X1  g412(.A(new_n534_), .B(G122), .ZN(G24));
  AOI21_X1  g413(.A(new_n519_), .B1(new_n472_), .B2(new_n471_), .ZN(new_n536_));
  NAND2_X1  g414(.A1(new_n511_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g415(.A(new_n537_), .B(G125), .ZN(G27));
  AOI21_X1  g416(.A(new_n522_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n539_));
  NOR2_X1   g417(.A1(new_n487_), .A2(new_n220_), .ZN(new_n540_));
  NAND3_X1  g418(.A1(new_n539_), .A2(new_n506_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g419(.A1(new_n541_), .A2(KEYINPUT40), .ZN(new_n542_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n543_));
  NAND4_X1  g421(.A1(new_n539_), .A2(new_n543_), .A3(new_n506_), .A4(new_n540_), .ZN(new_n544_));
  NAND2_X1  g422(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g423(.A(new_n545_), .B(new_n198_), .ZN(new_n546_));
  XNOR2_X1  g424(.A(new_n546_), .B(KEYINPUT41), .ZN(G33));
  NAND3_X1  g425(.A1(new_n539_), .A2(new_n484_), .A3(new_n540_), .ZN(new_n548_));
  XNOR2_X1  g426(.A(new_n548_), .B(G134), .ZN(G36));
  NAND3_X1  g427(.A1(new_n454_), .A2(new_n441_), .A3(new_n363_), .ZN(new_n550_));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n551_));
  NAND2_X1  g429(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g430(.A1(new_n454_), .A2(new_n441_), .A3(KEYINPUT42), .A4(new_n363_), .ZN(new_n553_));
  NAND3_X1  g431(.A1(new_n552_), .A2(new_n446_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g432(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g433(.A1(new_n540_), .A2(new_n469_), .ZN(new_n556_));
  NOR3_X1   g434(.A1(new_n398_), .A2(new_n390_), .A3(new_n388_), .ZN(new_n557_));
  NOR2_X1   g435(.A1(new_n422_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g436(.A(G469), .B1(new_n558_), .B2(G902), .ZN(new_n559_));
  AOI21_X1  g437(.A(new_n418_), .B1(new_n559_), .B2(new_n413_), .ZN(new_n560_));
  INV_X1    g438(.A(new_n483_), .ZN(new_n561_));
  NAND2_X1  g439(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g440(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g441(.A(KEYINPUT43), .B1(new_n555_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n565_));
  NOR4_X1   g443(.A1(new_n554_), .A2(new_n556_), .A3(new_n565_), .A4(new_n562_), .ZN(new_n566_));
  NOR2_X1   g444(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g445(.A(new_n567_), .B(G137), .Z(new_n568_));
  XNOR2_X1  g446(.A(new_n568_), .B(KEYINPUT44), .ZN(G39));
  NOR2_X1   g447(.A1(new_n521_), .A2(new_n446_), .ZN(new_n570_));
  NAND3_X1  g448(.A1(new_n506_), .A2(new_n560_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g449(.A(new_n540_), .ZN(new_n572_));
  NOR2_X1   g450(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g451(.A(new_n573_), .B(new_n144_), .ZN(new_n574_));
  XNOR2_X1  g452(.A(new_n574_), .B(KEYINPUT45), .ZN(G42));
  AND2_X1   g453(.A1(new_n545_), .A2(new_n548_), .ZN(new_n576_));
  AOI21_X1  g454(.A(new_n449_), .B1(new_n421_), .B2(new_n434_), .ZN(new_n577_));
  AOI21_X1  g455(.A(new_n460_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n578_));
  NAND2_X1  g456(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g457(.A(new_n579_), .ZN(new_n580_));
  AND3_X1   g458(.A1(new_n432_), .A2(KEYINPUT49), .A3(new_n561_), .ZN(new_n581_));
  AOI21_X1  g459(.A(KEYINPUT49), .B1(new_n432_), .B2(new_n561_), .ZN(new_n582_));
  NOR2_X1   g460(.A1(new_n442_), .A2(new_n455_), .ZN(new_n583_));
  XNOR2_X1  g461(.A(new_n583_), .B(KEYINPUT50), .ZN(new_n584_));
  AND3_X1   g462(.A1(new_n584_), .A2(new_n480_), .A3(new_n540_), .ZN(new_n585_));
  INV_X1    g463(.A(new_n498_), .ZN(new_n586_));
  NOR4_X1   g464(.A1(new_n586_), .A2(new_n510_), .A3(new_n469_), .A4(new_n491_), .ZN(new_n587_));
  OAI22_X1  g465(.A1(new_n581_), .A2(new_n582_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  AND4_X1   g466(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .A4(new_n534_), .ZN(new_n589_));
  NAND4_X1  g467(.A1(new_n432_), .A2(new_n473_), .A3(new_n506_), .A4(new_n540_), .ZN(new_n590_));
  NAND3_X1  g468(.A1(new_n589_), .A2(new_n485_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g469(.A1(new_n512_), .A2(new_n537_), .ZN(new_n592_));
  NOR2_X1   g470(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g471(.A1(new_n576_), .A2(new_n580_), .A3(new_n588_), .A4(new_n593_), .ZN(new_n594_));
  INV_X1    g472(.A(new_n594_), .ZN(new_n595_));
  AND2_X1   g473(.A1(new_n552_), .A2(new_n553_), .ZN(new_n596_));
  INV_X1    g474(.A(new_n278_), .ZN(new_n597_));
  AND3_X1   g475(.A1(new_n596_), .A2(new_n597_), .A3(new_n520_), .ZN(new_n598_));
  INV_X1    g476(.A(new_n448_), .ZN(new_n599_));
  NAND2_X1  g477(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g478(.A1(new_n600_), .A2(G952), .A3(new_n141_), .ZN(new_n601_));
  XNOR2_X1  g479(.A(new_n601_), .B(KEYINPUT47), .ZN(new_n602_));
  NAND4_X1  g480(.A1(new_n598_), .A2(new_n220_), .A3(new_n447_), .A4(new_n489_), .ZN(new_n603_));
  NAND3_X1  g481(.A1(new_n595_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g482(.A1(new_n531_), .A2(new_n418_), .ZN(new_n605_));
  NOR2_X1   g483(.A1(new_n605_), .A2(KEYINPUT48), .ZN(new_n606_));
  NOR2_X1   g484(.A1(new_n606_), .A2(new_n560_), .ZN(new_n607_));
  NAND2_X1  g485(.A1(new_n605_), .A2(KEYINPUT48), .ZN(new_n608_));
  AOI211_X1 g486(.A(new_n446_), .B(new_n165_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g487(.A(new_n597_), .B(new_n596_), .C1(new_n609_), .C2(new_n536_), .ZN(new_n610_));
  NAND2_X1  g488(.A1(new_n444_), .A2(KEYINPUT46), .ZN(new_n611_));
  OAI21_X1  g489(.A(new_n611_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n612_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n613_));
  NAND2_X1  g491(.A1(new_n443_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g492(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g493(.A(new_n586_), .B1(new_n612_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g494(.A1(new_n616_), .A2(new_n554_), .ZN(new_n617_));
  NAND4_X1  g495(.A1(new_n617_), .A2(new_n521_), .A3(new_n597_), .A4(new_n520_), .ZN(new_n618_));
  AOI21_X1  g496(.A(new_n572_), .B1(new_n610_), .B2(new_n618_), .ZN(new_n619_));
  OAI22_X1  g497(.A1(new_n604_), .A2(new_n619_), .B1(G952), .B2(G953), .ZN(new_n620_));
  NOR3_X1   g498(.A1(new_n498_), .A2(new_n165_), .A3(new_n500_), .ZN(new_n621_));
  AND3_X1   g499(.A1(new_n441_), .A2(new_n363_), .A3(new_n309_), .ZN(new_n622_));
  NAND4_X1  g500(.A1(new_n621_), .A2(new_n489_), .A3(new_n531_), .A4(new_n622_), .ZN(new_n623_));
  NAND2_X1  g501(.A1(new_n620_), .A2(new_n623_), .ZN(G75));
  NOR2_X1   g502(.A1(new_n141_), .A2(G952), .ZN(new_n625_));
  INV_X1    g503(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g504(.A1(new_n274_), .A2(new_n158_), .ZN(new_n627_));
  OR2_X1    g505(.A1(new_n262_), .A2(new_n265_), .ZN(new_n628_));
  NAND3_X1  g506(.A1(new_n628_), .A2(KEYINPUT51), .A3(new_n266_), .ZN(new_n629_));
  NAND3_X1  g507(.A1(new_n594_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g508(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g509(.A(new_n629_), .B1(new_n594_), .B2(new_n627_), .ZN(new_n632_));
  OAI21_X1  g510(.A(new_n626_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g511(.A(new_n633_), .B(KEYINPUT52), .ZN(G51));
  NOR2_X1   g512(.A1(new_n412_), .A2(new_n158_), .ZN(new_n635_));
  NAND4_X1  g513(.A1(new_n593_), .A2(new_n545_), .A3(new_n548_), .A4(new_n588_), .ZN(new_n636_));
  OAI211_X1 g514(.A(new_n558_), .B(new_n635_), .C1(new_n636_), .C2(new_n579_), .ZN(new_n637_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n638_));
  NAND2_X1  g516(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g517(.A1(new_n594_), .A2(KEYINPUT53), .A3(new_n558_), .A4(new_n635_), .ZN(new_n640_));
  NAND2_X1  g518(.A1(new_n594_), .A2(new_n635_), .ZN(new_n641_));
  AOI22_X1  g519(.A1(new_n639_), .A2(new_n640_), .B1(new_n641_), .B2(new_n411_), .ZN(new_n642_));
  OR3_X1    g520(.A1(new_n642_), .A2(KEYINPUT54), .A3(new_n625_), .ZN(new_n643_));
  OAI21_X1  g521(.A(KEYINPUT54), .B1(new_n642_), .B2(new_n625_), .ZN(new_n644_));
  NAND2_X1  g522(.A1(new_n643_), .A2(new_n644_), .ZN(G54));
  NAND3_X1  g523(.A1(new_n594_), .A2(G475), .A3(G902), .ZN(new_n646_));
  NOR2_X1   g524(.A1(new_n361_), .A2(new_n362_), .ZN(new_n647_));
  XNOR2_X1  g525(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  NOR2_X1   g526(.A1(new_n648_), .A2(new_n625_), .ZN(G60));
  NAND3_X1  g527(.A1(new_n594_), .A2(G478), .A3(G902), .ZN(new_n650_));
  XOR2_X1   g528(.A(new_n650_), .B(new_n349_), .Z(new_n651_));
  NOR2_X1   g529(.A1(new_n651_), .A2(new_n625_), .ZN(G63));
  INV_X1    g530(.A(new_n162_), .ZN(new_n653_));
  NOR2_X1   g531(.A1(new_n160_), .A2(new_n158_), .ZN(new_n654_));
  NAND3_X1  g532(.A1(new_n594_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g533(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g534(.A(new_n653_), .B1(new_n594_), .B2(new_n654_), .ZN(new_n657_));
  OAI21_X1  g535(.A(new_n626_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n659_));
  XNOR2_X1  g537(.A(new_n658_), .B(new_n659_), .ZN(G66));
  AOI21_X1  g538(.A(new_n137_), .B1(G224), .B2(G898), .ZN(new_n661_));
  INV_X1    g539(.A(new_n661_), .ZN(new_n662_));
  NAND4_X1  g540(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .A4(new_n534_), .ZN(new_n663_));
  NAND2_X1  g541(.A1(new_n663_), .A2(KEYINPUT56), .ZN(new_n664_));
  NAND2_X1  g542(.A1(new_n218_), .A2(new_n276_), .ZN(new_n665_));
  NOR2_X1   g543(.A1(new_n665_), .A2(new_n519_), .ZN(new_n666_));
  AOI22_X1  g544(.A1(new_n666_), .A2(new_n458_), .B1(new_n528_), .B2(new_n520_), .ZN(new_n667_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n668_));
  NAND4_X1  g546(.A1(new_n667_), .A2(new_n668_), .A3(new_n524_), .A4(new_n534_), .ZN(new_n669_));
  NAND2_X1  g547(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g548(.A1(new_n577_), .A2(new_n578_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n672_));
  NAND2_X1  g550(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g551(.A1(new_n577_), .A2(new_n578_), .A3(new_n670_), .A4(KEYINPUT57), .ZN(new_n674_));
  NAND3_X1  g552(.A1(new_n673_), .A2(new_n137_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g553(.A1(new_n675_), .A2(KEYINPUT58), .ZN(new_n676_));
  INV_X1    g554(.A(KEYINPUT58), .ZN(new_n677_));
  NAND4_X1  g555(.A1(new_n673_), .A2(new_n677_), .A3(new_n137_), .A4(new_n674_), .ZN(new_n678_));
  INV_X1    g556(.A(new_n141_), .ZN(new_n679_));
  AOI21_X1  g557(.A(new_n265_), .B1(new_n280_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g558(.A1(new_n676_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g559(.A(new_n680_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n682_));
  INV_X1    g560(.A(KEYINPUT59), .ZN(new_n683_));
  OAI21_X1  g561(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI211_X1 g562(.A(KEYINPUT59), .B(new_n680_), .C1(new_n676_), .C2(new_n678_), .ZN(new_n685_));
  OAI21_X1  g563(.A(new_n662_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g564(.A1(new_n680_), .A2(new_n662_), .ZN(new_n687_));
  XOR2_X1   g565(.A(new_n687_), .B(KEYINPUT60), .Z(new_n688_));
  NAND2_X1  g566(.A1(new_n686_), .A2(new_n688_), .ZN(G69));
  NOR2_X1   g567(.A1(new_n567_), .A2(new_n573_), .ZN(new_n690_));
  NAND3_X1  g568(.A1(new_n545_), .A2(new_n690_), .A3(new_n548_), .ZN(new_n691_));
  INV_X1    g569(.A(KEYINPUT61), .ZN(new_n692_));
  NAND2_X1  g570(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g571(.A1(new_n545_), .A2(new_n690_), .A3(KEYINPUT61), .A4(new_n548_), .ZN(new_n694_));
  NAND4_X1  g572(.A1(new_n523_), .A2(new_n561_), .A3(new_n490_), .A4(new_n560_), .ZN(new_n695_));
  AND4_X1   g573(.A1(new_n485_), .A2(new_n512_), .A3(new_n537_), .A4(new_n695_), .ZN(new_n696_));
  NAND3_X1  g574(.A1(new_n693_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g575(.A1(new_n697_), .A2(new_n137_), .ZN(new_n698_));
  XOR2_X1   g576(.A(new_n210_), .B(new_n148_), .Z(new_n699_));
  AOI21_X1  g577(.A(new_n699_), .B1(new_n481_), .B2(G953), .ZN(new_n700_));
  NAND2_X1  g578(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g579(.A(new_n141_), .B1(G227), .B2(G900), .ZN(new_n702_));
  NAND2_X1  g580(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g581(.A1(new_n700_), .A2(new_n679_), .ZN(new_n704_));
  NAND3_X1  g582(.A1(new_n611_), .A2(new_n456_), .A3(new_n614_), .ZN(new_n705_));
  NAND4_X1  g583(.A1(new_n432_), .A2(new_n218_), .A3(new_n561_), .A4(new_n705_), .ZN(new_n706_));
  AOI21_X1  g584(.A(new_n572_), .B1(new_n706_), .B2(new_n571_), .ZN(new_n707_));
  INV_X1    g585(.A(new_n537_), .ZN(new_n708_));
  NOR4_X1   g586(.A1(new_n504_), .A2(new_n707_), .A3(new_n708_), .A4(new_n567_), .ZN(new_n709_));
  NAND3_X1  g587(.A1(new_n709_), .A2(new_n485_), .A3(new_n512_), .ZN(new_n710_));
  AOI22_X1  g588(.A1(new_n698_), .A2(new_n700_), .B1(new_n704_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g589(.A(new_n703_), .B1(new_n711_), .B2(new_n702_), .ZN(G72));
  NOR2_X1   g590(.A1(new_n166_), .A2(new_n158_), .ZN(new_n713_));
  XNOR2_X1  g591(.A(new_n713_), .B(KEYINPUT62), .ZN(new_n714_));
  NAND4_X1  g592(.A1(new_n709_), .A2(new_n485_), .A3(new_n512_), .A4(new_n589_), .ZN(new_n715_));
  OAI21_X1  g593(.A(new_n714_), .B1(new_n715_), .B2(new_n579_), .ZN(new_n716_));
  OAI211_X1 g594(.A(new_n495_), .B(new_n713_), .C1(new_n636_), .C2(new_n579_), .ZN(new_n717_));
  INV_X1    g595(.A(KEYINPUT63), .ZN(new_n718_));
  NAND2_X1  g596(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND4_X1  g597(.A1(new_n594_), .A2(KEYINPUT63), .A3(new_n495_), .A4(new_n713_), .ZN(new_n720_));
  AOI22_X1  g598(.A1(new_n494_), .A2(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g599(.A(new_n181_), .ZN(new_n722_));
  OAI21_X1  g600(.A(new_n626_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  AND2_X1   g601(.A1(new_n673_), .A2(new_n674_), .ZN(new_n724_));
  OAI21_X1  g602(.A(new_n714_), .B1(new_n697_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g603(.A1(new_n725_), .A2(new_n495_), .ZN(new_n726_));
  NAND3_X1  g604(.A1(new_n594_), .A2(new_n494_), .A3(new_n713_), .ZN(new_n727_));
  AOI21_X1  g605(.A(new_n181_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g606(.A1(new_n723_), .A2(new_n728_), .ZN(G57));
endmodule


