//Secret key is'0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_c1355" written by ABC on Wed Nov 16 09:08:33 2022

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat,
    G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203_));
  AND2_X1   g002(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NOR4_X1   g007(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT65), .A4(G190gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT63), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT62), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT63), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT62), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n202_), .B1(new_n210_), .B2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n220_), .A2(new_n221_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT64), .B(G183gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT65), .B1(new_n225_), .B2(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n206_), .A2(new_n203_), .A3(new_n207_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n228_), .A3(KEYINPUT66), .ZN(new_n229_));
  INV_X1    g028(.A(new_n221_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n215_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT60), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT59), .B(G176gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n234_), .B1(new_n235_), .B2(new_n212_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n213_), .A2(KEYINPUT59), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT59), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G176gat), .ZN(new_n239_));
  AND4_X1   g038(.A1(new_n234_), .A2(new_n237_), .A3(new_n239_), .A4(new_n212_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n233_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT61), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n239_), .A3(new_n212_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT60), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n235_), .A2(new_n234_), .A3(new_n212_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT61), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n233_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n223_), .A2(new_n229_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  INV_X1    g049(.A(G120gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G113gat), .ZN(new_n252_));
  INV_X1    g051(.A(G113gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G120gat), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256_));
  INV_X1    g055(.A(G127gat), .ZN(new_n257_));
  INV_X1    g056(.A(G134gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(G127gat), .B2(G134gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G127gat), .A2(G134gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT3), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n256_), .B(new_n259_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT2), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n255_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(KEYINPUT3), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n260_), .A2(G127gat), .A3(G134gat), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n267_), .A2(new_n268_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n252_), .A2(new_n254_), .A3(new_n265_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n256_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n250_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n256_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n259_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT2), .B1(new_n269_), .B2(new_n256_), .ZN(new_n276_));
  OAI211_X1 g075(.A(KEYINPUT12), .B(new_n275_), .C1(new_n276_), .C2(new_n255_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n249_), .A2(new_n272_), .A3(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n224_), .A2(new_n228_), .A3(KEYINPUT66), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT66), .B1(new_n224_), .B2(new_n228_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n247_), .B1(new_n246_), .B2(new_n233_), .ZN(new_n281_));
  AOI211_X1 g080(.A(KEYINPUT61), .B(new_n232_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n282_));
  OAI22_X1  g081(.A1(new_n279_), .A2(new_n280_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n272_), .A2(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n278_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G227gat), .A2(G233gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n278_), .A2(new_n285_), .A3(new_n288_), .A4(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT73), .Z(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(KEYINPUT75), .A3(new_n298_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT76), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT76), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n306_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G1gat), .B(G29gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT0), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n275_), .B1(new_n276_), .B2(new_n255_), .ZN(new_n314_));
  INV_X1    g113(.A(G155gat), .ZN(new_n315_));
  INV_X1    g114(.A(G162gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT7), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G155gat), .A3(G162gat), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n317_), .A2(KEYINPUT8), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT8), .B1(new_n317_), .B2(new_n319_), .ZN(new_n321_));
  OAI22_X1  g120(.A1(new_n320_), .A2(new_n321_), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT6), .B(G141gat), .ZN(new_n323_));
  INV_X1    g122(.A(G148gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT5), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT11), .ZN(new_n330_));
  OR2_X1    g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n317_), .A2(new_n319_), .B1(new_n331_), .B2(new_n326_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT10), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT9), .B(G155gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n316_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n315_), .A2(KEYINPUT9), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G155gat), .ZN(new_n338_));
  AND4_X1   g137(.A1(new_n333_), .A2(new_n336_), .A3(new_n338_), .A4(new_n316_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n330_), .B(new_n332_), .C1(new_n335_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n338_), .A3(new_n316_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT10), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n336_), .A2(new_n338_), .A3(new_n333_), .A4(new_n316_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n330_), .B1(new_n345_), .B2(new_n332_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n314_), .B(new_n329_), .C1(new_n341_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT14), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n332_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT11), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n340_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT14), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n329_), .A4(new_n314_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n348_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT13), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n351_), .A2(new_n340_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(new_n284_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n329_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(KEYINPUT13), .A3(new_n272_), .A4(new_n277_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(KEYINPUT15), .A3(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n357_), .A2(new_n314_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n347_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n349_), .B(KEYINPUT1), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT15), .B1(new_n355_), .B2(new_n361_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n313_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n355_), .A2(new_n361_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT15), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(new_n312_), .A3(new_n366_), .A4(new_n362_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G197gat), .ZN(new_n378_));
  INV_X1    g177(.A(G204gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT53), .A2(G197gat), .A3(G204gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT53), .B1(G197gat), .B2(G204gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G211gat), .A2(G218gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT55), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT54), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT54), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(G211gat), .A3(G218gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n384_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G218gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT56), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT56), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G218gat), .ZN(new_n396_));
  INV_X1    g195(.A(G211gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT57), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT57), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n394_), .A2(new_n396_), .A3(new_n400_), .A4(new_n397_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(new_n384_), .A3(new_n391_), .A4(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT58), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT53), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n381_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(KEYINPUT57), .A2(new_n398_), .B1(new_n408_), .B2(new_n380_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n401_), .A2(new_n391_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(KEYINPUT58), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n392_), .B1(new_n404_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G228gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT71), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  AOI211_X1 g215(.A(new_n392_), .B(new_n414_), .C1(new_n404_), .C2(new_n411_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n359_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n392_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n402_), .A2(new_n403_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT58), .B1(new_n409_), .B2(new_n410_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n414_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n412_), .A2(new_n415_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n357_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(new_n425_), .A3(KEYINPUT70), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT72), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G22gat), .B(G50gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n418_), .A2(new_n425_), .A3(KEYINPUT70), .A4(new_n430_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n427_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n377_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n428_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n376_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(new_n249_), .B2(new_n412_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n283_), .A2(new_n422_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT68), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n283_), .A2(new_n422_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n249_), .A2(new_n412_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT68), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .A4(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n283_), .B2(new_n422_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n249_), .A2(KEYINPUT67), .A3(new_n412_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n444_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n440_), .B(KEYINPUT52), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G8gat), .B(G36gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT50), .B(KEYINPUT51), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n448_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n308_), .A2(new_n375_), .A3(new_n439_), .A4(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT77), .ZN(new_n469_));
  INV_X1    g268(.A(new_n308_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n434_), .A2(new_n438_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n467_), .A3(new_n375_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n462_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n455_), .A2(new_n473_), .A3(new_n461_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n374_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n365_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n363_), .A2(KEYINPUT80), .A3(new_n347_), .A4(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n348_), .A2(new_n354_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n349_), .B1(new_n482_), .B2(new_n361_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n479_), .B(new_n481_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n313_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n462_), .A2(new_n464_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n373_), .A3(new_n488_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n477_), .A2(new_n489_), .B1(new_n438_), .B2(new_n434_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n472_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n477_), .A2(new_n489_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n493_), .A2(new_n491_), .A3(new_n439_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n470_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(KEYINPUT82), .B(new_n470_), .C1(new_n492_), .C2(new_n494_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n469_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT17), .B1(G85gat), .B2(G92gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G85gat), .ZN(new_n505_));
  INV_X1    g304(.A(G92gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT22), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OR3_X1    g306(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT22), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT19), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n509_), .B(new_n511_), .C1(G99gat), .C2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n504_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n502_), .A2(new_n503_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT18), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n514_), .A2(new_n516_), .B1(G85gat), .B2(G92gat), .ZN(new_n517_));
  INV_X1    g316(.A(G99gat), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n511_), .A2(KEYINPUT20), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n510_), .B(KEYINPUT19), .Z(new_n521_));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n517_), .A2(KEYINPUT21), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT21), .B1(new_n517_), .B2(new_n524_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n512_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G29gat), .B(G36gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(G50gat), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n533_), .A2(G43gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT33), .B(G43gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(G50gat), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n532_), .A2(KEYINPUT34), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n530_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT34), .B(new_n538_), .C1(new_n532_), .C2(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(KEYINPUT43), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(KEYINPUT43), .ZN(new_n542_));
  OAI211_X1 g341(.A(KEYINPUT28), .B(new_n512_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n529_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n540_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n527_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G134gat), .B(G162gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT83), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT84), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT85), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n545_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n548_), .B(new_n555_), .C1(new_n556_), .C2(KEYINPUT86), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n556_), .A2(KEYINPUT86), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT87), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n544_), .A2(new_n547_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n545_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT86), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n548_), .A2(new_n555_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n556_), .A2(KEYINPUT86), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n559_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n554_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n562_), .B2(new_n548_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n499_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT23), .Z(new_n576_));
  NOR2_X1   g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G57gat), .A2(G64gat), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT26), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  INV_X1    g381(.A(G57gat), .ZN(new_n583_));
  INV_X1    g382(.A(G64gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n578_), .B1(new_n581_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n576_), .A2(KEYINPUT24), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n576_), .A2(KEYINPUT24), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n577_), .B(KEYINPUT25), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n579_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n587_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n527_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G230gat), .ZN(new_n595_));
  INV_X1    g394(.A(G233gat), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n529_), .A2(new_n543_), .A3(new_n593_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT29), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT29), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n529_), .A2(new_n602_), .A3(new_n543_), .A4(new_n593_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n599_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n527_), .A2(new_n593_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT27), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT27), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n527_), .A2(new_n607_), .A3(new_n593_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n598_), .B1(new_n609_), .B2(new_n594_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n604_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G120gat), .B(G148gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n611_), .A2(KEYINPUT30), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n604_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n610_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n616_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n615_), .B1(new_n604_), .B2(new_n610_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(KEYINPUT30), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT39), .B(G22gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT38), .B(G15gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G1gat), .A2(G8gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(KEYINPUT37), .A2(G1gat), .A3(G8gat), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n631_), .B(new_n632_), .C1(G1gat), .C2(G8gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G15gat), .A2(G22gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(G15gat), .A2(G22gat), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n634_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n639_), .B2(new_n634_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G1gat), .Z(new_n642_));
  OAI211_X1 g441(.A(new_n641_), .B(new_n629_), .C1(G8gat), .C2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n635_), .A2(new_n636_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n637_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n625_), .B1(new_n645_), .B2(new_n540_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n637_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n546_), .A2(KEYINPUT41), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n540_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(KEYINPUT42), .A3(new_n540_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(G229gat), .A2(G233gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n645_), .A2(KEYINPUT44), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n647_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n541_), .A2(new_n658_), .A3(new_n542_), .A4(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n655_), .A3(new_n650_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G169gat), .B(G197gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT31), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n667_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n657_), .A2(new_n662_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n624_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n593_), .A2(new_n647_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT48), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n658_), .A2(new_n660_), .A3(new_n593_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(G231gat), .A2(G233gat), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT47), .Z(new_n678_));
  OAI211_X1 g477(.A(new_n675_), .B(new_n676_), .C1(KEYINPUT49), .C2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT49), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(G127gat), .B(G155gat), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT46), .ZN(new_n684_));
  XNOR2_X1  g483(.A(G183gat), .B(G211gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n681_), .B(new_n686_), .Z(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n574_), .A2(new_n673_), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G1gat), .B1(new_n689_), .B2(new_n375_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n469_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n493_), .A2(new_n439_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT81), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n490_), .A2(new_n491_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n472_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT82), .B1(new_n695_), .B2(new_n470_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n498_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n691_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT89), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT89), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n499_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(new_n671_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT90), .B1(new_n569_), .B2(new_n572_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT90), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n705_), .B(new_n571_), .C1(new_n559_), .C2(new_n568_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n624_), .A3(new_n687_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n703_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n374_), .B(KEYINPUT88), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(new_n642_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n690_), .B1(new_n710_), .B2(new_n713_), .ZN(G1324gat));
  INV_X1    g513(.A(G8gat), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n689_), .A2(new_n715_), .A3(new_n467_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n467_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n703_), .A2(new_n717_), .A3(new_n709_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n715_), .ZN(G1325gat));
  AND4_X1   g518(.A1(new_n308_), .A2(new_n703_), .A3(new_n627_), .A4(new_n709_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT91), .ZN(new_n721_));
  OAI21_X1  g520(.A(G15gat), .B1(new_n689_), .B2(new_n470_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1326gat));
  AND4_X1   g522(.A1(new_n471_), .A2(new_n703_), .A3(new_n626_), .A4(new_n709_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT93), .ZN(new_n725_));
  OAI21_X1  g524(.A(G22gat), .B1(new_n689_), .B2(new_n439_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT92), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1327gat));
  NAND2_X1  g527(.A1(new_n687_), .A2(new_n573_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n624_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n703_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G29gat), .B1(new_n732_), .B2(new_n711_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT94), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n698_), .A2(new_n734_), .A3(new_n708_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT94), .B1(new_n499_), .B2(new_n707_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n688_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n673_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n374_), .A2(G29gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n733_), .B1(new_n738_), .B2(new_n739_), .ZN(G1328gat));
  AOI21_X1  g539(.A(G36gat), .B1(new_n732_), .B2(new_n717_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n717_), .A2(G36gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n738_), .B2(new_n742_), .ZN(G1329gat));
  NAND4_X1  g542(.A1(new_n703_), .A2(new_n535_), .A3(new_n308_), .A4(new_n730_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n308_), .A3(new_n673_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n745_), .A2(KEYINPUT95), .A3(G43gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT95), .B1(new_n745_), .B2(G43gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT96), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(G1330gat));
  OAI21_X1  g549(.A(new_n533_), .B1(new_n731_), .B2(new_n439_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n738_), .A2(G50gat), .A3(new_n471_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT97), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT97), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n755_), .A3(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1331gat));
  AND2_X1   g556(.A1(new_n624_), .A2(KEYINPUT98), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n624_), .A2(KEYINPUT98), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n687_), .A2(new_n671_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR4_X1   g561(.A1(new_n499_), .A2(new_n573_), .A3(new_n760_), .A4(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n374_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G57gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT99), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n762_), .A2(new_n708_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n702_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT100), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n702_), .A2(KEYINPUT100), .A3(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n760_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n711_), .A2(new_n583_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n767_), .B(new_n768_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n760_), .B(new_n777_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT101), .B1(new_n779_), .B2(new_n766_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1332gat));
  AOI21_X1  g580(.A(new_n584_), .B1(new_n763_), .B2(new_n717_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n760_), .A2(new_n467_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n584_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n782_), .B1(new_n774_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT102), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(G1333gat));
  INV_X1    g587(.A(G71gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n763_), .B2(new_n308_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT103), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n308_), .A2(new_n789_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n776_), .B2(new_n792_), .ZN(G1334gat));
  INV_X1    g592(.A(G78gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n763_), .B2(new_n471_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT104), .Z(new_n796_));
  NAND2_X1  g595(.A1(new_n471_), .A2(new_n794_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n776_), .B2(new_n797_), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n760_), .A2(new_n671_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n737_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n374_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G85gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n729_), .A2(new_n671_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n699_), .A2(new_n701_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT105), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n699_), .A2(new_n701_), .A3(new_n806_), .A4(new_n803_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n760_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n505_), .A3(new_n711_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n802_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1336gat));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n807_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n506_), .A3(new_n783_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n800_), .A2(new_n717_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n506_), .ZN(G1337gat));
  NAND3_X1  g615(.A1(new_n808_), .A2(new_n518_), .A3(new_n308_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n800_), .A2(new_n308_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n518_), .ZN(G1338gat));
  NOR2_X1   g618(.A1(new_n439_), .A2(G106gat), .ZN(new_n820_));
  AND4_X1   g619(.A1(KEYINPUT108), .A2(new_n813_), .A3(new_n775_), .A4(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT108), .B1(new_n808_), .B2(new_n820_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT107), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n735_), .A2(new_n736_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(new_n471_), .A3(new_n687_), .A4(new_n799_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n825_), .B2(G106gat), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n825_), .A2(new_n823_), .A3(G106gat), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n821_), .A2(new_n822_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT109), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n830_));
  OAI221_X1 g629(.A(new_n830_), .B1(new_n826_), .B2(new_n827_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1339gat));
  AOI21_X1  g631(.A(new_n655_), .B1(new_n661_), .B2(new_n650_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n834_));
  OAI22_X1  g633(.A1(new_n833_), .A2(new_n834_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT112), .B(new_n655_), .C1(new_n661_), .C2(new_n650_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n666_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n670_), .A2(KEYINPUT111), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n657_), .A2(new_n839_), .A3(new_n662_), .A4(new_n669_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n620_), .A2(new_n837_), .A3(new_n838_), .A4(new_n840_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n604_), .A2(KEYINPUT110), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n604_), .A2(KEYINPUT110), .ZN(new_n843_));
  INV_X1    g642(.A(new_n594_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n842_), .B(new_n843_), .C1(new_n598_), .C2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n841_), .B1(new_n615_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n837_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n617_), .A3(new_n622_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n604_), .A2(KEYINPUT110), .B1(new_n845_), .B2(new_n598_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n843_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n615_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n671_), .A3(new_n620_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n573_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n848_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI211_X1 g656(.A(KEYINPUT113), .B(new_n573_), .C1(new_n850_), .C2(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n687_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n761_), .A2(new_n623_), .A3(new_n707_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n471_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n861_), .A2(KEYINPUT114), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n712_), .A2(new_n717_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(KEYINPUT114), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n862_), .A2(new_n308_), .A3(new_n863_), .A4(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(new_n253_), .A3(new_n672_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n859_), .A2(new_n860_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT115), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n859_), .A2(new_n869_), .A3(new_n860_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n712_), .ZN(new_n872_));
  AND4_X1   g671(.A1(new_n308_), .A2(new_n872_), .A3(new_n439_), .A4(new_n467_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n671_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n866_), .B1(new_n874_), .B2(new_n253_), .ZN(G1340gat));
  XOR2_X1   g674(.A(KEYINPUT116), .B(G120gat), .Z(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n775_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G120gat), .B1(new_n865_), .B2(new_n623_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(KEYINPUT117), .A3(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1341gat));
  NOR3_X1   g682(.A1(new_n865_), .A2(new_n257_), .A3(new_n687_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n873_), .A2(new_n688_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n257_), .ZN(G1342gat));
  NAND3_X1  g685(.A1(new_n873_), .A2(new_n258_), .A3(new_n573_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G134gat), .B1(new_n865_), .B2(new_n707_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n888_), .A2(KEYINPUT118), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n888_), .A2(KEYINPUT118), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n887_), .B1(new_n890_), .B2(new_n891_), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n308_), .A2(new_n439_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n867_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n863_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895_), .B2(new_n672_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT119), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n872_), .A2(new_n467_), .A3(new_n893_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n671_), .A2(new_n323_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1344gat));
  OAI21_X1  g699(.A(new_n324_), .B1(new_n898_), .B2(new_n760_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n894_), .A2(G148gat), .A3(new_n624_), .A4(new_n863_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n895_), .B2(new_n687_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n688_), .A2(new_n334_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n898_), .B2(new_n907_), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n895_), .B2(new_n707_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT121), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n573_), .A2(new_n316_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n898_), .A2(new_n911_), .ZN(new_n912_));
  MUX2_X1   g711(.A(new_n910_), .B(KEYINPUT121), .S(new_n912_), .Z(G1347gat));
  NOR4_X1   g712(.A1(new_n871_), .A2(new_n374_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n467_), .A2(new_n672_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n914_), .A2(new_n212_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n467_), .A2(new_n374_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n862_), .A2(new_n308_), .A3(new_n864_), .A4(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G169gat), .B1(new_n920_), .B2(new_n672_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n917_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n918_), .A2(new_n921_), .A3(new_n922_), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n914_), .A2(new_n235_), .A3(new_n783_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G176gat), .B1(new_n920_), .B2(new_n623_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1349gat));
  NAND4_X1  g725(.A1(new_n914_), .A2(new_n206_), .A3(new_n717_), .A4(new_n688_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G183gat), .B1(new_n920_), .B2(new_n687_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1350gat));
  NAND4_X1  g728(.A1(new_n914_), .A2(new_n207_), .A3(new_n573_), .A4(new_n717_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G190gat), .B1(new_n920_), .B2(new_n707_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1351gat));
  NAND2_X1  g731(.A1(new_n894_), .A2(new_n919_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933_), .B2(new_n672_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n859_), .A2(new_n869_), .A3(new_n860_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n869_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n937_), .A2(KEYINPUT123), .A3(new_n375_), .A4(new_n893_), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n868_), .A2(new_n375_), .A3(new_n870_), .A4(new_n893_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n915_), .A2(new_n378_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n934_), .B1(new_n943_), .B2(new_n944_), .ZN(G1352gat));
  OAI21_X1  g744(.A(G204gat), .B1(new_n933_), .B2(new_n623_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  OAI211_X1 g747(.A(KEYINPUT124), .B(G204gat), .C1(new_n933_), .C2(new_n623_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n783_), .A2(new_n379_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(KEYINPUT125), .B1(new_n942_), .B2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954_));
  AOI211_X1 g753(.A(new_n954_), .B(new_n951_), .C1(new_n938_), .C2(new_n941_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n950_), .B1(new_n953_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  OAI211_X1 g757(.A(KEYINPUT126), .B(new_n950_), .C1(new_n953_), .C2(new_n955_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1353gat));
  NOR3_X1   g759(.A1(new_n687_), .A2(G211gat), .A3(new_n467_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n942_), .A2(new_n961_), .ZN(new_n962_));
  OR2_X1    g761(.A1(new_n962_), .A2(KEYINPUT127), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(KEYINPUT127), .ZN(new_n964_));
  OAI21_X1  g763(.A(G211gat), .B1(new_n933_), .B2(new_n687_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n933_), .B2(new_n707_), .ZN(new_n967_));
  NAND4_X1  g766(.A1(new_n573_), .A2(new_n394_), .A3(new_n396_), .A4(new_n717_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n967_), .B1(new_n943_), .B2(new_n968_), .ZN(G1355gat));
endmodule


