//Secret key is'1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_c3540" written by ABC on Wed Nov 16 09:45:49 2022

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G13, G20, G33, G41, G45, G50, G58, G68,
    G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150,
    G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244,
    G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326,
    G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G13, G20, G33, G41, G45,
    G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201_, new_n202_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1222_, new_n1223_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201_));
  INV_X1    g0001(.A(G77), .ZN(new_n202_));
  AND2_X1   g0002(.A1(new_n201_), .A2(new_n202_), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205_));
  NOR2_X1   g0005(.A1(new_n205_), .A2(G13), .ZN(new_n206_));
  OAI211_X1 g0006(.A(new_n206_), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207_));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208_));
  XNOR2_X1  g0008(.A(new_n208_), .B(KEYINPUT3), .ZN(new_n209_));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210_));
  NAND2_X1  g0010(.A1(new_n210_), .A2(G20), .ZN(new_n211_));
  OAI21_X1  g0011(.A(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g0012(.A(G68), .ZN(new_n213_));
  INV_X1    g0013(.A(G238), .ZN(new_n214_));
  INV_X1    g0014(.A(G87), .ZN(new_n215_));
  INV_X1    g0015(.A(G250), .ZN(new_n216_));
  OAI22_X1  g0016(.A1(new_n213_), .A2(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g0017(.A1(G77), .A2(G244), .ZN(new_n218_));
  INV_X1    g0018(.A(G107), .ZN(new_n219_));
  INV_X1    g0019(.A(G264), .ZN(new_n220_));
  OAI21_X1  g0020(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222_));
  INV_X1    g0022(.A(G58), .ZN(new_n223_));
  INV_X1    g0023(.A(G232), .ZN(new_n224_));
  OAI21_X1  g0024(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NOR3_X1   g0025(.A1(new_n217_), .A2(new_n221_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g0026(.A(G50), .ZN(new_n227_));
  XOR2_X1   g0027(.A(KEYINPUT0), .B(G226), .Z(new_n228_));
  XNOR2_X1  g0028(.A(KEYINPUT1), .B(G97), .ZN(new_n229_));
  INV_X1    g0029(.A(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G257), .ZN(new_n231_));
  OAI221_X1 g0031(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g0032(.A(new_n212_), .B1(new_n232_), .B2(new_n205_), .ZN(G361));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234_));
  XNOR2_X1  g0034(.A(new_n234_), .B(KEYINPUT4), .ZN(new_n235_));
  XNOR2_X1  g0035(.A(new_n235_), .B(KEYINPUT5), .ZN(new_n236_));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237_));
  XNOR2_X1  g0037(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239_));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240_));
  XNOR2_X1  g0040(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g0041(.A(new_n238_), .B(new_n241_), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243_));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244_));
  XNOR2_X1  g0044(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246_));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247_));
  XNOR2_X1  g0047(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g0048(.A(new_n245_), .B(new_n248_), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT30), .ZN(new_n250_));
  NOR2_X1   g0050(.A1(G33), .A2(G1698), .ZN(new_n251_));
  AOI22_X1  g0051(.A1(new_n251_), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n252_));
  INV_X1    g0052(.A(G33), .ZN(new_n253_));
  NAND2_X1  g0053(.A1(new_n253_), .A2(G1698), .ZN(new_n254_));
  OAI21_X1  g0054(.A(new_n252_), .B1(new_n228_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g0055(.A1(G33), .A2(G41), .ZN(new_n256_));
  NAND2_X1  g0056(.A1(G1), .A2(G13), .ZN(new_n257_));
  NOR2_X1   g0057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g0058(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g0059(.A(KEYINPUT8), .B1(new_n256_), .B2(new_n257_), .ZN(new_n260_));
  INV_X1    g0060(.A(KEYINPUT8), .ZN(new_n261_));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262_));
  NAND3_X1  g0062(.A1(new_n210_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g0063(.A(G1), .ZN(new_n264_));
  OAI21_X1  g0064(.A(new_n264_), .B1(G41), .B2(G45), .ZN(new_n265_));
  NAND4_X1  g0065(.A1(new_n260_), .A2(new_n263_), .A3(G232), .A4(new_n265_), .ZN(new_n266_));
  OAI211_X1 g0066(.A(new_n264_), .B(G274), .C1(G41), .C2(G45), .ZN(new_n267_));
  NAND3_X1  g0067(.A1(new_n259_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g0068(.A1(new_n268_), .A2(G169), .ZN(new_n269_));
  NAND2_X1  g0069(.A1(new_n269_), .A2(KEYINPUT31), .ZN(new_n270_));
  INV_X1    g0070(.A(KEYINPUT31), .ZN(new_n271_));
  NAND3_X1  g0071(.A1(new_n268_), .A2(new_n271_), .A3(G169), .ZN(new_n272_));
  INV_X1    g0072(.A(G179), .ZN(new_n273_));
  OR2_X1    g0073(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g0074(.A1(new_n270_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g0075(.A1(new_n257_), .A2(KEYINPUT10), .ZN(new_n276_));
  INV_X1    g0076(.A(KEYINPUT10), .ZN(new_n277_));
  NAND3_X1  g0077(.A1(new_n277_), .A2(G1), .A3(G13), .ZN(new_n278_));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279_));
  AND3_X1   g0079(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g0080(.A(G20), .ZN(new_n281_));
  NAND3_X1  g0081(.A1(new_n281_), .A2(G33), .A3(G68), .ZN(new_n282_));
  INV_X1    g0082(.A(KEYINPUT28), .ZN(new_n283_));
  XNOR2_X1  g0083(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g0084(.A(G58), .B(G68), .ZN(new_n285_));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286_));
  AOI22_X1  g0086(.A1(new_n285_), .A2(G20), .B1(G159), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g0087(.A(new_n280_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g0088(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g0089(.A(KEYINPUT29), .ZN(new_n290_));
  NAND3_X1  g0090(.A1(new_n264_), .A2(G13), .A3(G20), .ZN(new_n291_));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292_));
  NAND2_X1  g0092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g0093(.A1(new_n264_), .A2(KEYINPUT9), .A3(G13), .A4(G20), .ZN(new_n294_));
  NAND2_X1  g0094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g0095(.A1(new_n281_), .A2(G1), .ZN(new_n296_));
  INV_X1    g0096(.A(new_n296_), .ZN(new_n297_));
  NAND4_X1  g0097(.A1(new_n295_), .A2(new_n280_), .A3(G58), .A4(new_n297_), .ZN(new_n298_));
  NAND3_X1  g0098(.A1(new_n289_), .A2(new_n290_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g0099(.A(new_n298_), .ZN(new_n300_));
  OAI21_X1  g0100(.A(KEYINPUT29), .B1(new_n300_), .B2(new_n288_), .ZN(new_n301_));
  NAND2_X1  g0101(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g0102(.A1(new_n293_), .A2(new_n294_), .ZN(new_n303_));
  NAND2_X1  g0103(.A1(new_n303_), .A2(new_n223_), .ZN(new_n304_));
  NAND2_X1  g0104(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g0105(.A1(new_n275_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g0106(.A1(new_n268_), .A2(G200), .ZN(new_n307_));
  INV_X1    g0107(.A(G190), .ZN(new_n308_));
  NOR2_X1   g0108(.A1(new_n268_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g0109(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g0110(.A1(new_n299_), .A2(new_n301_), .B1(new_n223_), .B2(new_n303_), .ZN(new_n311_));
  NAND2_X1  g0111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g0112(.A(new_n250_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g0113(.A(KEYINPUT30), .B1(new_n310_), .B2(new_n311_), .ZN(new_n314_));
  NOR2_X1   g0114(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g0115(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g0116(.A1(new_n295_), .A2(new_n280_), .ZN(new_n317_));
  INV_X1    g0117(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g0118(.A1(new_n318_), .A2(G50), .A3(new_n297_), .ZN(new_n319_));
  NAND2_X1  g0119(.A1(new_n281_), .A2(G33), .ZN(new_n320_));
  INV_X1    g0120(.A(new_n320_), .ZN(new_n321_));
  AOI22_X1  g0121(.A1(new_n321_), .A2(G58), .B1(new_n286_), .B2(G150), .ZN(new_n322_));
  OAI21_X1  g0122(.A(new_n322_), .B1(new_n281_), .B2(new_n201_), .ZN(new_n323_));
  NAND3_X1  g0123(.A1(new_n276_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n324_));
  AOI22_X1  g0124(.A1(new_n323_), .A2(new_n324_), .B1(new_n303_), .B2(new_n227_), .ZN(new_n325_));
  AND2_X1   g0125(.A1(new_n260_), .A2(new_n263_), .ZN(new_n326_));
  NAND3_X1  g0126(.A1(new_n326_), .A2(G226), .A3(new_n265_), .ZN(new_n327_));
  INV_X1    g0127(.A(G1698), .ZN(new_n328_));
  NOR2_X1   g0128(.A1(new_n328_), .A2(G33), .ZN(new_n329_));
  AOI22_X1  g0129(.A1(new_n329_), .A2(G223), .B1(G33), .B2(G77), .ZN(new_n330_));
  INV_X1    g0130(.A(G222), .ZN(new_n331_));
  INV_X1    g0131(.A(new_n251_), .ZN(new_n332_));
  OAI21_X1  g0132(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g0133(.A1(new_n333_), .A2(new_n258_), .ZN(new_n334_));
  NAND3_X1  g0134(.A1(new_n327_), .A2(new_n334_), .A3(new_n267_), .ZN(new_n335_));
  OAI211_X1 g0135(.A(new_n319_), .B(new_n325_), .C1(new_n335_), .C2(new_n308_), .ZN(new_n336_));
  AND2_X1   g0136(.A1(new_n335_), .A2(G200), .ZN(new_n337_));
  NOR2_X1   g0137(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OR2_X1    g0138(.A1(new_n338_), .A2(KEYINPUT14), .ZN(new_n339_));
  NAND2_X1  g0139(.A1(new_n338_), .A2(KEYINPUT14), .ZN(new_n340_));
  INV_X1    g0140(.A(G169), .ZN(new_n341_));
  NAND2_X1  g0141(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g0142(.A1(new_n325_), .A2(new_n319_), .ZN(new_n343_));
  OAI211_X1 g0143(.A(new_n342_), .B(new_n343_), .C1(G179), .C2(new_n335_), .ZN(new_n344_));
  NAND3_X1  g0144(.A1(new_n339_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g0145(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g0146(.A1(new_n228_), .A2(new_n332_), .ZN(new_n347_));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348_));
  OR2_X1    g0148(.A1(new_n348_), .A2(KEYINPUT17), .ZN(new_n349_));
  NAND2_X1  g0149(.A1(new_n348_), .A2(KEYINPUT17), .ZN(new_n350_));
  OAI211_X1 g0150(.A(new_n349_), .B(new_n350_), .C1(new_n224_), .C2(new_n254_), .ZN(new_n351_));
  OAI21_X1  g0151(.A(new_n258_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g0152(.A1(new_n326_), .A2(G238), .A3(new_n265_), .ZN(new_n353_));
  NAND4_X1  g0153(.A1(new_n352_), .A2(new_n353_), .A3(G190), .A4(new_n267_), .ZN(new_n354_));
  AOI21_X1  g0154(.A(G20), .B1(G33), .B2(G77), .ZN(new_n355_));
  NAND2_X1  g0155(.A1(new_n253_), .A2(G50), .ZN(new_n356_));
  AOI22_X1  g0156(.A1(new_n355_), .A2(new_n356_), .B1(G20), .B2(G68), .ZN(new_n357_));
  NAND2_X1  g0157(.A1(new_n357_), .A2(new_n324_), .ZN(new_n358_));
  XOR2_X1   g0158(.A(new_n358_), .B(KEYINPUT15), .Z(new_n359_));
  NAND3_X1  g0159(.A1(new_n303_), .A2(KEYINPUT16), .A3(new_n213_), .ZN(new_n360_));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361_));
  OAI21_X1  g0161(.A(new_n361_), .B1(new_n295_), .B2(G68), .ZN(new_n362_));
  NAND2_X1  g0162(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g0163(.A1(new_n318_), .A2(G68), .A3(new_n297_), .ZN(new_n364_));
  NAND4_X1  g0164(.A1(new_n354_), .A2(new_n359_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366_));
  NAND3_X1  g0166(.A1(new_n352_), .A2(new_n353_), .A3(new_n267_), .ZN(new_n367_));
  AOI21_X1  g0167(.A(new_n366_), .B1(new_n367_), .B2(G200), .ZN(new_n368_));
  INV_X1    g0168(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g0169(.A1(new_n367_), .A2(new_n366_), .A3(G200), .ZN(new_n370_));
  AOI21_X1  g0170(.A(new_n365_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g0171(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n372_));
  NAND4_X1  g0172(.A1(new_n352_), .A2(new_n353_), .A3(new_n273_), .A4(new_n267_), .ZN(new_n373_));
  NAND2_X1  g0173(.A1(new_n367_), .A2(new_n341_), .ZN(new_n374_));
  NAND3_X1  g0174(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g0175(.A(new_n375_), .ZN(new_n376_));
  OAI21_X1  g0176(.A(KEYINPUT19), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g0177(.A(new_n372_), .ZN(new_n378_));
  INV_X1    g0178(.A(new_n370_), .ZN(new_n379_));
  OAI211_X1 g0179(.A(new_n378_), .B(new_n354_), .C1(new_n379_), .C2(new_n368_), .ZN(new_n380_));
  INV_X1    g0180(.A(KEYINPUT19), .ZN(new_n381_));
  NAND3_X1  g0181(.A1(new_n380_), .A2(new_n381_), .A3(new_n375_), .ZN(new_n382_));
  NAND2_X1  g0182(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g0183(.A1(new_n346_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g0184(.A1(new_n303_), .A2(new_n202_), .ZN(new_n385_));
  NAND3_X1  g0185(.A1(new_n318_), .A2(G77), .A3(new_n297_), .ZN(new_n386_));
  XNOR2_X1  g0186(.A(KEYINPUT20), .B(G87), .ZN(new_n387_));
  NAND3_X1  g0187(.A1(new_n387_), .A2(KEYINPUT21), .A3(new_n321_), .ZN(new_n388_));
  AOI22_X1  g0188(.A1(new_n286_), .A2(G58), .B1(G20), .B2(G77), .ZN(new_n389_));
  NAND2_X1  g0189(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g0190(.A(KEYINPUT21), .B1(new_n387_), .B2(new_n321_), .ZN(new_n391_));
  OAI21_X1  g0191(.A(new_n324_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g0192(.A(KEYINPUT22), .ZN(new_n393_));
  AND2_X1   g0193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g0194(.A(KEYINPUT22), .B(new_n324_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n395_));
  INV_X1    g0195(.A(new_n395_), .ZN(new_n396_));
  OAI211_X1 g0196(.A(new_n385_), .B(new_n386_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g0197(.A(KEYINPUT11), .ZN(new_n398_));
  NOR2_X1   g0198(.A1(new_n398_), .A2(G107), .ZN(new_n399_));
  NOR2_X1   g0199(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n400_));
  OAI21_X1  g0200(.A(G33), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AOI22_X1  g0201(.A1(new_n329_), .A2(G238), .B1(new_n251_), .B2(G232), .ZN(new_n402_));
  INV_X1    g0202(.A(KEYINPUT23), .ZN(new_n403_));
  NAND3_X1  g0203(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g0204(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n405_));
  NAND2_X1  g0205(.A1(new_n398_), .A2(G107), .ZN(new_n406_));
  AOI21_X1  g0206(.A(new_n253_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g0207(.A1(new_n253_), .A2(new_n328_), .A3(G232), .ZN(new_n408_));
  NAND3_X1  g0208(.A1(new_n253_), .A2(G238), .A3(G1698), .ZN(new_n409_));
  NAND2_X1  g0209(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g0210(.A(KEYINPUT23), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g0211(.A1(new_n404_), .A2(new_n411_), .A3(new_n258_), .ZN(new_n412_));
  NAND4_X1  g0212(.A1(new_n260_), .A2(new_n263_), .A3(G244), .A4(new_n265_), .ZN(new_n413_));
  AND2_X1   g0213(.A1(new_n413_), .A2(new_n267_), .ZN(new_n414_));
  NAND2_X1  g0214(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g0215(.A(KEYINPUT24), .ZN(new_n416_));
  NAND2_X1  g0216(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g0217(.A1(new_n412_), .A2(new_n414_), .A3(KEYINPUT24), .ZN(new_n418_));
  AND3_X1   g0218(.A1(new_n417_), .A2(G169), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g0219(.A(KEYINPUT25), .ZN(new_n420_));
  OAI21_X1  g0220(.A(new_n420_), .B1(new_n415_), .B2(new_n273_), .ZN(new_n421_));
  NAND4_X1  g0221(.A1(new_n412_), .A2(new_n414_), .A3(KEYINPUT25), .A4(G179), .ZN(new_n422_));
  NAND2_X1  g0222(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g0223(.A(KEYINPUT26), .B(new_n397_), .C1(new_n419_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g0224(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g0225(.A1(new_n417_), .A2(G169), .A3(new_n418_), .ZN(new_n426_));
  NAND3_X1  g0226(.A1(new_n426_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n427_));
  AOI21_X1  g0227(.A(KEYINPUT26), .B1(new_n427_), .B2(new_n397_), .ZN(new_n428_));
  NOR2_X1   g0228(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g0229(.A(new_n397_), .ZN(new_n430_));
  NAND3_X1  g0230(.A1(new_n417_), .A2(G200), .A3(new_n418_), .ZN(new_n431_));
  OAI211_X1 g0231(.A(new_n430_), .B(new_n431_), .C1(new_n308_), .C2(new_n415_), .ZN(new_n432_));
  NAND2_X1  g0232(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g0233(.A(KEYINPUT27), .ZN(new_n434_));
  OR3_X1    g0234(.A1(new_n384_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  OAI21_X1  g0235(.A(new_n434_), .B1(new_n384_), .B2(new_n433_), .ZN(new_n436_));
  AOI21_X1  g0236(.A(new_n316_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g0237(.A1(new_n264_), .A2(G33), .ZN(new_n438_));
  NAND3_X1  g0238(.A1(new_n318_), .A2(new_n387_), .A3(new_n438_), .ZN(new_n439_));
  OAI211_X1 g0239(.A(new_n348_), .B(new_n281_), .C1(G33), .C2(new_n213_), .ZN(new_n440_));
  INV_X1    g0240(.A(G97), .ZN(new_n441_));
  NAND3_X1  g0241(.A1(new_n215_), .A2(new_n441_), .A3(new_n219_), .ZN(new_n442_));
  OAI211_X1 g0242(.A(new_n324_), .B(new_n440_), .C1(new_n281_), .C2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g0243(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g0244(.A1(new_n444_), .A2(KEYINPUT35), .ZN(new_n445_));
  INV_X1    g0245(.A(new_n387_), .ZN(new_n446_));
  NAND2_X1  g0246(.A1(new_n303_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g0247(.A(KEYINPUT35), .ZN(new_n448_));
  NAND3_X1  g0248(.A1(new_n439_), .A2(new_n448_), .A3(new_n443_), .ZN(new_n449_));
  NAND3_X1  g0249(.A1(new_n445_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g0250(.A(G45), .ZN(new_n451_));
  NOR2_X1   g0251(.A1(new_n451_), .A2(G1), .ZN(new_n452_));
  NOR2_X1   g0252(.A1(new_n452_), .A2(new_n216_), .ZN(new_n453_));
  NAND3_X1  g0253(.A1(new_n253_), .A2(G244), .A3(G1698), .ZN(new_n454_));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455_));
  OAI211_X1 g0255(.A(new_n454_), .B(new_n455_), .C1(new_n332_), .C2(new_n214_), .ZN(new_n456_));
  AOI22_X1  g0256(.A1(new_n326_), .A2(new_n453_), .B1(new_n258_), .B2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g0257(.A1(new_n260_), .A2(new_n263_), .A3(G274), .A4(new_n452_), .ZN(new_n458_));
  INV_X1    g0258(.A(KEYINPUT32), .ZN(new_n459_));
  AND2_X1   g0259(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g0260(.A1(new_n458_), .A2(new_n459_), .ZN(new_n461_));
  OAI21_X1  g0261(.A(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g0262(.A1(new_n462_), .A2(KEYINPUT33), .ZN(new_n463_));
  XNOR2_X1  g0263(.A(new_n458_), .B(new_n459_), .ZN(new_n464_));
  INV_X1    g0264(.A(KEYINPUT33), .ZN(new_n465_));
  NAND3_X1  g0265(.A1(new_n464_), .A2(new_n465_), .A3(new_n457_), .ZN(new_n466_));
  AND3_X1   g0266(.A1(new_n463_), .A2(G169), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g0267(.A(KEYINPUT34), .ZN(new_n468_));
  OAI21_X1  g0268(.A(new_n468_), .B1(new_n462_), .B2(new_n273_), .ZN(new_n469_));
  NAND4_X1  g0269(.A1(new_n464_), .A2(KEYINPUT34), .A3(G179), .A4(new_n457_), .ZN(new_n470_));
  NAND2_X1  g0270(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g0271(.A(new_n450_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g0272(.A(G41), .ZN(new_n473_));
  NAND3_X1  g0273(.A1(new_n264_), .A2(new_n473_), .A3(G45), .ZN(new_n474_));
  NAND4_X1  g0274(.A1(new_n260_), .A2(new_n263_), .A3(G257), .A4(new_n474_), .ZN(new_n475_));
  NAND3_X1  g0275(.A1(new_n260_), .A2(G274), .A3(new_n263_), .ZN(new_n476_));
  NAND3_X1  g0276(.A1(new_n452_), .A2(KEYINPUT7), .A3(new_n473_), .ZN(new_n477_));
  INV_X1    g0277(.A(KEYINPUT7), .ZN(new_n478_));
  NAND2_X1  g0278(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g0279(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g0280(.A(new_n475_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g0281(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g0282(.A1(new_n253_), .A2(new_n328_), .A3(G244), .ZN(new_n483_));
  NAND3_X1  g0283(.A1(new_n253_), .A2(G250), .A3(G1698), .ZN(new_n484_));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485_));
  NAND3_X1  g0285(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AND3_X1   g0286(.A1(new_n486_), .A2(KEYINPUT6), .A3(new_n258_), .ZN(new_n487_));
  AOI21_X1  g0287(.A(KEYINPUT6), .B1(new_n486_), .B2(new_n258_), .ZN(new_n488_));
  NOR2_X1   g0288(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g0289(.A1(new_n482_), .A2(G190), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g0290(.A1(new_n486_), .A2(new_n258_), .ZN(new_n491_));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g0292(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g0293(.A1(new_n486_), .A2(KEYINPUT6), .A3(new_n258_), .ZN(new_n494_));
  NAND2_X1  g0294(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g0295(.A(G200), .B1(new_n495_), .B2(new_n481_), .ZN(new_n496_));
  NAND3_X1  g0296(.A1(new_n230_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n497_));
  NAND2_X1  g0297(.A1(new_n438_), .A2(G97), .ZN(new_n498_));
  OAI21_X1  g0298(.A(new_n497_), .B1(new_n317_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g0299(.A1(new_n405_), .A2(new_n406_), .A3(G97), .ZN(new_n500_));
  OAI211_X1 g0300(.A(new_n500_), .B(G20), .C1(new_n219_), .C2(new_n229_), .ZN(new_n501_));
  AOI22_X1  g0301(.A1(new_n321_), .A2(G107), .B1(new_n286_), .B2(G77), .ZN(new_n502_));
  AOI21_X1  g0302(.A(new_n280_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g0303(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g0304(.A1(new_n490_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g0305(.A(KEYINPUT12), .ZN(new_n506_));
  NAND2_X1  g0306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g0307(.A1(new_n490_), .A2(new_n496_), .A3(new_n504_), .A4(KEYINPUT12), .ZN(new_n508_));
  INV_X1    g0308(.A(new_n499_), .ZN(new_n509_));
  INV_X1    g0309(.A(KEYINPUT13), .ZN(new_n510_));
  AND2_X1   g0310(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g0311(.A1(new_n503_), .A2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g0312(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g0313(.A(G169), .B1(new_n482_), .B2(new_n489_), .ZN(new_n514_));
  NOR3_X1   g0314(.A1(new_n495_), .A2(new_n481_), .A3(G179), .ZN(new_n515_));
  NOR2_X1   g0315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g0316(.A1(new_n507_), .A2(new_n508_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g0317(.A1(new_n462_), .A2(new_n308_), .ZN(new_n518_));
  NAND3_X1  g0318(.A1(new_n318_), .A2(G87), .A3(new_n438_), .ZN(new_n519_));
  NAND3_X1  g0319(.A1(new_n519_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n520_));
  NOR2_X1   g0320(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g0321(.A(G200), .ZN(new_n522_));
  NAND2_X1  g0322(.A1(new_n463_), .A2(new_n466_), .ZN(new_n523_));
  OAI21_X1  g0323(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g0324(.A1(new_n472_), .A2(new_n517_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g0325(.A1(new_n253_), .A2(new_n328_), .A3(G250), .ZN(new_n526_));
  NAND3_X1  g0326(.A1(new_n253_), .A2(G257), .A3(G1698), .ZN(new_n527_));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528_));
  NAND3_X1  g0328(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g0329(.A(KEYINPUT40), .ZN(new_n530_));
  AND3_X1   g0330(.A1(new_n529_), .A2(new_n530_), .A3(new_n258_), .ZN(new_n531_));
  AOI21_X1  g0331(.A(new_n530_), .B1(new_n529_), .B2(new_n258_), .ZN(new_n532_));
  OAI22_X1  g0332(.A1(new_n531_), .A2(new_n532_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n533_));
  NAND4_X1  g0333(.A1(new_n260_), .A2(new_n263_), .A3(G264), .A4(new_n474_), .ZN(new_n534_));
  NAND2_X1  g0334(.A1(new_n534_), .A2(G179), .ZN(new_n535_));
  OAI21_X1  g0335(.A(KEYINPUT41), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g0336(.A(new_n534_), .ZN(new_n537_));
  OAI21_X1  g0337(.A(G169), .B1(new_n533_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g0338(.A(new_n532_), .ZN(new_n539_));
  NAND3_X1  g0339(.A1(new_n529_), .A2(new_n530_), .A3(new_n258_), .ZN(new_n540_));
  NAND2_X1  g0340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g0341(.A(new_n535_), .ZN(new_n542_));
  AND2_X1   g0342(.A1(new_n477_), .A2(new_n479_), .ZN(new_n543_));
  NAND3_X1  g0343(.A1(new_n543_), .A2(new_n326_), .A3(G274), .ZN(new_n544_));
  INV_X1    g0344(.A(KEYINPUT41), .ZN(new_n545_));
  NAND4_X1  g0345(.A1(new_n541_), .A2(new_n542_), .A3(new_n544_), .A4(new_n545_), .ZN(new_n546_));
  NAND3_X1  g0346(.A1(new_n536_), .A2(new_n538_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g0347(.A1(new_n405_), .A2(new_n406_), .ZN(new_n548_));
  AOI21_X1  g0348(.A(G20), .B1(new_n293_), .B2(new_n294_), .ZN(new_n549_));
  NOR3_X1   g0349(.A1(new_n318_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g0350(.A1(new_n253_), .A2(G87), .ZN(new_n551_));
  AOI21_X1  g0351(.A(G20), .B1(new_n551_), .B2(new_n455_), .ZN(new_n552_));
  NAND2_X1  g0352(.A1(new_n324_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g0353(.A1(new_n438_), .A2(G107), .ZN(new_n554_));
  OAI21_X1  g0354(.A(new_n553_), .B1(new_n317_), .B2(new_n554_), .ZN(new_n555_));
  OR2_X1    g0355(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g0356(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g0357(.A(KEYINPUT42), .ZN(new_n558_));
  NAND2_X1  g0358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g0359(.A1(new_n547_), .A2(new_n556_), .A3(KEYINPUT42), .ZN(new_n560_));
  NOR2_X1   g0360(.A1(new_n550_), .A2(new_n555_), .ZN(new_n561_));
  NAND3_X1  g0361(.A1(new_n541_), .A2(new_n544_), .A3(new_n534_), .ZN(new_n562_));
  NAND2_X1  g0362(.A1(new_n562_), .A2(G200), .ZN(new_n563_));
  OAI211_X1 g0363(.A(new_n561_), .B(new_n563_), .C1(new_n562_), .C2(new_n308_), .ZN(new_n564_));
  NAND3_X1  g0364(.A1(new_n559_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g0365(.A1(new_n525_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g0366(.A(KEYINPUT37), .ZN(new_n567_));
  INV_X1    g0367(.A(KEYINPUT36), .ZN(new_n568_));
  INV_X1    g0368(.A(G283), .ZN(new_n569_));
  OAI21_X1  g0369(.A(new_n568_), .B1(new_n320_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g0370(.A1(KEYINPUT1), .A2(G97), .ZN(new_n571_));
  NOR2_X1   g0371(.A1(KEYINPUT1), .A2(G97), .ZN(new_n572_));
  OAI21_X1  g0372(.A(new_n286_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g0373(.A1(G20), .A2(G116), .ZN(new_n574_));
  NAND4_X1  g0374(.A1(new_n281_), .A2(KEYINPUT36), .A3(G33), .A4(G283), .ZN(new_n575_));
  NAND4_X1  g0375(.A1(new_n570_), .A2(new_n573_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NAND2_X1  g0376(.A1(new_n576_), .A2(new_n324_), .ZN(new_n577_));
  NAND4_X1  g0377(.A1(new_n295_), .A2(new_n280_), .A3(G116), .A4(new_n438_), .ZN(new_n578_));
  INV_X1    g0378(.A(G116), .ZN(new_n579_));
  NAND2_X1  g0379(.A1(new_n303_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g0380(.A1(new_n577_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g0381(.A(new_n581_), .ZN(new_n582_));
  NAND4_X1  g0382(.A1(new_n260_), .A2(new_n263_), .A3(G270), .A4(new_n474_), .ZN(new_n583_));
  NOR2_X1   g0383(.A1(new_n231_), .A2(new_n332_), .ZN(new_n584_));
  INV_X1    g0384(.A(G303), .ZN(new_n585_));
  OAI22_X1  g0385(.A1(new_n254_), .A2(new_n220_), .B1(new_n253_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g0386(.A(new_n258_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g0387(.A1(new_n544_), .A2(G179), .A3(new_n583_), .A4(new_n587_), .ZN(new_n588_));
  OAI21_X1  g0388(.A(new_n567_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g0389(.A1(new_n476_), .A2(new_n480_), .ZN(new_n590_));
  INV_X1    g0390(.A(new_n258_), .ZN(new_n591_));
  INV_X1    g0391(.A(G257), .ZN(new_n592_));
  AND2_X1   g0392(.A1(new_n592_), .A2(KEYINPUT2), .ZN(new_n593_));
  NOR2_X1   g0393(.A1(new_n592_), .A2(KEYINPUT2), .ZN(new_n594_));
  OAI21_X1  g0394(.A(new_n251_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  AOI22_X1  g0395(.A1(new_n329_), .A2(G264), .B1(G33), .B2(G303), .ZN(new_n596_));
  AOI21_X1  g0396(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g0397(.A(new_n583_), .ZN(new_n598_));
  NOR3_X1   g0398(.A1(new_n590_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND4_X1  g0399(.A1(new_n599_), .A2(KEYINPUT37), .A3(new_n581_), .A4(G179), .ZN(new_n600_));
  NAND2_X1  g0400(.A1(new_n589_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g0401(.A(KEYINPUT38), .ZN(new_n602_));
  NAND3_X1  g0402(.A1(new_n544_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n603_));
  NAND3_X1  g0403(.A1(new_n603_), .A2(new_n581_), .A3(G169), .ZN(new_n604_));
  AND3_X1   g0404(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g0405(.A(new_n602_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n606_));
  OAI21_X1  g0406(.A(new_n582_), .B1(new_n603_), .B2(new_n308_), .ZN(new_n607_));
  INV_X1    g0407(.A(KEYINPUT39), .ZN(new_n608_));
  OAI21_X1  g0408(.A(new_n608_), .B1(new_n599_), .B2(new_n522_), .ZN(new_n609_));
  NAND3_X1  g0409(.A1(new_n603_), .A2(KEYINPUT39), .A3(G200), .ZN(new_n610_));
  AOI21_X1  g0410(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g0411(.A1(new_n605_), .A2(new_n606_), .A3(new_n611_), .ZN(new_n612_));
  AND3_X1   g0412(.A1(new_n437_), .A2(new_n566_), .A3(new_n612_), .ZN(G372));
  NAND2_X1  g0413(.A1(new_n339_), .A2(new_n340_), .ZN(new_n614_));
  OAI21_X1  g0414(.A(new_n344_), .B1(new_n614_), .B2(new_n306_), .ZN(new_n615_));
  NOR3_X1   g0415(.A1(new_n384_), .A2(new_n316_), .A3(new_n429_), .ZN(new_n616_));
  XOR2_X1   g0416(.A(new_n375_), .B(KEYINPUT43), .Z(new_n617_));
  NOR2_X1   g0417(.A1(new_n617_), .A2(new_n345_), .ZN(new_n618_));
  AOI211_X1 g0418(.A(new_n615_), .B(new_n616_), .C1(new_n315_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g0419(.A(new_n437_), .ZN(new_n620_));
  AND2_X1   g0420(.A1(new_n516_), .A2(new_n513_), .ZN(new_n621_));
  NAND2_X1  g0421(.A1(new_n524_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g0422(.A1(new_n622_), .A2(new_n472_), .ZN(new_n623_));
  AND3_X1   g0423(.A1(new_n472_), .A2(new_n517_), .A3(new_n524_), .ZN(new_n624_));
  NAND2_X1  g0424(.A1(new_n559_), .A2(new_n560_), .ZN(new_n625_));
  AOI21_X1  g0425(.A(new_n623_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g0426(.A(new_n565_), .ZN(new_n627_));
  NAND2_X1  g0427(.A1(new_n601_), .A2(new_n604_), .ZN(new_n628_));
  NAND3_X1  g0428(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g0429(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g0430(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g0431(.A(new_n619_), .B1(new_n620_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g0432(.A(new_n632_), .B(KEYINPUT44), .Z(G369));
  NOR2_X1   g0433(.A1(new_n605_), .A2(new_n606_), .ZN(new_n634_));
  INV_X1    g0434(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g0435(.A(G13), .ZN(new_n636_));
  INV_X1    g0436(.A(G213), .ZN(new_n637_));
  NOR4_X1   g0437(.A1(new_n636_), .A2(new_n637_), .A3(G1), .A4(G20), .ZN(new_n638_));
  INV_X1    g0438(.A(new_n638_), .ZN(new_n639_));
  INV_X1    g0439(.A(G343), .ZN(new_n640_));
  NOR2_X1   g0440(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g0441(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g0442(.A1(new_n582_), .A2(new_n642_), .ZN(new_n643_));
  MUX2_X1   g0443(.A(new_n612_), .B(new_n635_), .S(new_n643_), .Z(new_n644_));
  INV_X1    g0444(.A(KEYINPUT45), .ZN(new_n645_));
  NAND3_X1  g0445(.A1(new_n556_), .A2(new_n645_), .A3(new_n641_), .ZN(new_n646_));
  OAI21_X1  g0446(.A(KEYINPUT45), .B1(new_n561_), .B2(new_n642_), .ZN(new_n647_));
  NAND2_X1  g0447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OR2_X1    g0448(.A1(new_n648_), .A2(KEYINPUT46), .ZN(new_n649_));
  NAND2_X1  g0449(.A1(new_n648_), .A2(KEYINPUT46), .ZN(new_n650_));
  NAND2_X1  g0450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g0451(.A1(new_n651_), .A2(new_n565_), .ZN(new_n652_));
  NAND3_X1  g0452(.A1(new_n627_), .A2(new_n650_), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g0453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g0454(.A(KEYINPUT47), .B(G330), .Z(new_n655_));
  INV_X1    g0455(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g0456(.A1(new_n644_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g0457(.A(new_n634_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n658_));
  NOR2_X1   g0458(.A1(new_n658_), .A2(new_n625_), .ZN(new_n659_));
  OAI21_X1  g0459(.A(new_n657_), .B1(new_n659_), .B2(new_n641_), .ZN(G399));
  INV_X1    g0460(.A(KEYINPUT48), .ZN(new_n661_));
  INV_X1    g0461(.A(new_n206_), .ZN(new_n662_));
  OAI21_X1  g0462(.A(new_n661_), .B1(new_n662_), .B2(G41), .ZN(new_n663_));
  NAND3_X1  g0463(.A1(new_n206_), .A2(KEYINPUT48), .A3(new_n473_), .ZN(new_n664_));
  NAND2_X1  g0464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NOR3_X1   g0465(.A1(new_n665_), .A2(KEYINPUT49), .A3(new_n264_), .ZN(new_n666_));
  NOR3_X1   g0466(.A1(new_n666_), .A2(G116), .A3(new_n442_), .ZN(new_n667_));
  OAI21_X1  g0467(.A(KEYINPUT49), .B1(new_n665_), .B2(new_n264_), .ZN(new_n668_));
  INV_X1    g0468(.A(new_n209_), .ZN(new_n669_));
  AOI22_X1  g0469(.A1(new_n667_), .A2(new_n668_), .B1(new_n669_), .B2(new_n665_), .ZN(new_n670_));
  INV_X1    g0470(.A(KEYINPUT50), .ZN(new_n671_));
  NAND3_X1  g0471(.A1(new_n630_), .A2(new_n671_), .A3(new_n642_), .ZN(new_n672_));
  INV_X1    g0472(.A(new_n628_), .ZN(new_n673_));
  NOR3_X1   g0473(.A1(new_n525_), .A2(new_n565_), .A3(new_n673_), .ZN(new_n674_));
  OAI211_X1 g0474(.A(new_n469_), .B(new_n470_), .C1(new_n523_), .C2(new_n341_), .ZN(new_n675_));
  AOI22_X1  g0475(.A1(new_n524_), .A2(new_n621_), .B1(new_n675_), .B2(new_n450_), .ZN(new_n676_));
  INV_X1    g0476(.A(new_n560_), .ZN(new_n677_));
  AOI21_X1  g0477(.A(KEYINPUT42), .B1(new_n547_), .B2(new_n556_), .ZN(new_n678_));
  NOR2_X1   g0478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g0479(.A(new_n676_), .B1(new_n525_), .B2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g0480(.A(new_n642_), .B1(new_n674_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g0481(.A1(new_n681_), .A2(KEYINPUT50), .ZN(new_n682_));
  NAND2_X1  g0482(.A1(new_n672_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g0483(.A1(new_n624_), .A2(new_n612_), .A3(new_n627_), .A4(new_n642_), .ZN(new_n684_));
  INV_X1    g0484(.A(KEYINPUT51), .ZN(new_n685_));
  NAND2_X1  g0485(.A1(new_n482_), .A2(new_n489_), .ZN(new_n686_));
  NOR3_X1   g0486(.A1(new_n562_), .A2(new_n686_), .A3(new_n588_), .ZN(new_n687_));
  NAND2_X1  g0487(.A1(new_n687_), .A2(new_n523_), .ZN(new_n688_));
  NAND4_X1  g0488(.A1(new_n686_), .A2(new_n562_), .A3(new_n273_), .A4(new_n603_), .ZN(new_n689_));
  OAI21_X1  g0489(.A(new_n688_), .B1(new_n689_), .B2(new_n523_), .ZN(new_n690_));
  AOI21_X1  g0490(.A(new_n685_), .B1(new_n690_), .B2(new_n641_), .ZN(new_n691_));
  NAND2_X1  g0491(.A1(new_n684_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g0492(.A1(new_n566_), .A2(new_n685_), .A3(new_n612_), .A4(new_n642_), .ZN(new_n693_));
  NAND2_X1  g0493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g0494(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g0495(.A(new_n683_), .B1(G330), .B2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g0496(.A(new_n670_), .B1(new_n696_), .B2(G1), .ZN(G364));
  XNOR2_X1  g0497(.A(new_n644_), .B(G330), .ZN(new_n698_));
  XNOR2_X1  g0498(.A(new_n698_), .B(KEYINPUT52), .ZN(new_n699_));
  NAND2_X1  g0499(.A1(new_n699_), .A2(new_n665_), .ZN(new_n700_));
  XOR2_X1   g0500(.A(new_n700_), .B(KEYINPUT53), .Z(new_n701_));
  NOR2_X1   g0501(.A1(new_n636_), .A2(G20), .ZN(new_n702_));
  AOI21_X1  g0502(.A(new_n264_), .B1(new_n702_), .B2(G45), .ZN(new_n703_));
  XOR2_X1   g0503(.A(new_n703_), .B(KEYINPUT54), .Z(new_n704_));
  NAND2_X1  g0504(.A1(new_n699_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g0505(.A(new_n257_), .B1(G20), .B2(new_n341_), .ZN(new_n706_));
  OR2_X1    g0506(.A1(new_n706_), .A2(KEYINPUT60), .ZN(new_n707_));
  NAND2_X1  g0507(.A1(new_n706_), .A2(KEYINPUT60), .ZN(new_n708_));
  NAND2_X1  g0508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g0509(.A(new_n709_), .ZN(new_n710_));
  NOR3_X1   g0510(.A1(new_n281_), .A2(new_n273_), .A3(new_n308_), .ZN(new_n711_));
  INV_X1    g0511(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g0512(.A1(KEYINPUT56), .A2(G200), .ZN(new_n713_));
  INV_X1    g0513(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g0514(.A1(KEYINPUT56), .A2(G200), .ZN(new_n715_));
  NOR2_X1   g0515(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g0516(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g0517(.A1(new_n712_), .A2(G200), .ZN(new_n718_));
  AOI22_X1  g0518(.A1(G50), .A2(new_n717_), .B1(new_n718_), .B2(G58), .ZN(new_n719_));
  NOR2_X1   g0519(.A1(new_n281_), .A2(G190), .ZN(new_n720_));
  INV_X1    g0520(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g0521(.A1(new_n721_), .A2(new_n273_), .ZN(new_n722_));
  INV_X1    g0522(.A(new_n716_), .ZN(new_n723_));
  NAND2_X1  g0523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g0524(.A1(new_n722_), .A2(new_n716_), .ZN(new_n725_));
  OAI221_X1 g0525(.A(new_n719_), .B1(new_n213_), .B2(new_n724_), .C1(new_n202_), .C2(new_n725_), .ZN(new_n726_));
  XOR2_X1   g0526(.A(new_n726_), .B(KEYINPUT57), .Z(new_n727_));
  NOR3_X1   g0527(.A1(new_n716_), .A2(new_n721_), .A3(G179), .ZN(new_n728_));
  NAND2_X1  g0528(.A1(new_n728_), .A2(G107), .ZN(new_n729_));
  NOR2_X1   g0529(.A1(new_n281_), .A2(new_n308_), .ZN(new_n730_));
  NAND3_X1  g0530(.A1(new_n723_), .A2(new_n273_), .A3(new_n730_), .ZN(new_n731_));
  NOR2_X1   g0531(.A1(new_n731_), .A2(new_n215_), .ZN(new_n732_));
  NOR2_X1   g0532(.A1(new_n732_), .A2(G33), .ZN(new_n733_));
  OAI21_X1  g0533(.A(G20), .B1(G179), .B2(G200), .ZN(new_n734_));
  INV_X1    g0534(.A(KEYINPUT55), .ZN(new_n735_));
  XNOR2_X1  g0535(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  NOR2_X1   g0536(.A1(new_n736_), .A2(new_n720_), .ZN(new_n737_));
  INV_X1    g0537(.A(new_n737_), .ZN(new_n738_));
  NOR2_X1   g0538(.A1(new_n738_), .A2(new_n230_), .ZN(new_n739_));
  NOR2_X1   g0539(.A1(new_n736_), .A2(new_n721_), .ZN(new_n740_));
  AOI21_X1  g0540(.A(new_n739_), .B1(G159), .B2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g0541(.A1(new_n727_), .A2(new_n729_), .A3(new_n733_), .A4(new_n741_), .ZN(new_n742_));
  INV_X1    g0542(.A(new_n728_), .ZN(new_n743_));
  INV_X1    g0543(.A(G322), .ZN(new_n744_));
  INV_X1    g0544(.A(new_n718_), .ZN(new_n745_));
  OAI221_X1 g0545(.A(G33), .B1(new_n743_), .B2(new_n569_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n746_));
  INV_X1    g0546(.A(new_n731_), .ZN(new_n747_));
  AOI21_X1  g0547(.A(new_n746_), .B1(G303), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g0548(.A1(new_n740_), .A2(G329), .ZN(new_n749_));
  XNOR2_X1  g0549(.A(new_n749_), .B(KEYINPUT59), .ZN(new_n750_));
  NAND2_X1  g0550(.A1(new_n737_), .A2(G294), .ZN(new_n751_));
  INV_X1    g0551(.A(new_n717_), .ZN(new_n752_));
  INV_X1    g0552(.A(G326), .ZN(new_n753_));
  INV_X1    g0553(.A(G317), .ZN(new_n754_));
  OAI22_X1  g0554(.A1(new_n752_), .A2(new_n753_), .B1(new_n754_), .B2(new_n724_), .ZN(new_n755_));
  INV_X1    g0555(.A(new_n725_), .ZN(new_n756_));
  XNOR2_X1  g0556(.A(KEYINPUT58), .B(G311), .ZN(new_n757_));
  AOI21_X1  g0557(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g0558(.A1(new_n748_), .A2(new_n750_), .A3(new_n751_), .A4(new_n758_), .ZN(new_n759_));
  AOI21_X1  g0559(.A(new_n710_), .B1(new_n742_), .B2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761_));
  XOR2_X1   g0561(.A(new_n761_), .B(KEYINPUT62), .Z(new_n762_));
  NOR2_X1   g0562(.A1(new_n762_), .A2(G20), .ZN(new_n763_));
  INV_X1    g0563(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g0564(.A1(new_n764_), .A2(new_n710_), .ZN(new_n765_));
  NOR2_X1   g0565(.A1(new_n662_), .A2(new_n253_), .ZN(new_n766_));
  INV_X1    g0566(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g0567(.A(new_n767_), .B1(new_n669_), .B2(new_n451_), .ZN(new_n768_));
  OAI21_X1  g0568(.A(new_n768_), .B1(new_n248_), .B2(new_n451_), .ZN(new_n769_));
  XOR2_X1   g0569(.A(new_n769_), .B(KEYINPUT61), .Z(new_n770_));
  NOR2_X1   g0570(.A1(new_n662_), .A2(G33), .ZN(new_n771_));
  AOI22_X1  g0571(.A1(new_n771_), .A2(G355), .B1(new_n579_), .B2(new_n662_), .ZN(new_n772_));
  AOI21_X1  g0572(.A(new_n765_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g0573(.A1(new_n704_), .A2(new_n665_), .ZN(new_n774_));
  INV_X1    g0574(.A(new_n774_), .ZN(new_n775_));
  NOR3_X1   g0575(.A1(new_n760_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g0576(.A(new_n776_), .B1(new_n644_), .B2(new_n764_), .ZN(new_n777_));
  NAND3_X1  g0577(.A1(new_n701_), .A2(new_n705_), .A3(new_n777_), .ZN(G396));
  NAND2_X1  g0578(.A1(new_n397_), .A2(new_n641_), .ZN(new_n779_));
  INV_X1    g0579(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g0580(.A(new_n780_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n781_));
  OAI21_X1  g0581(.A(new_n397_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n782_));
  INV_X1    g0582(.A(KEYINPUT26), .ZN(new_n783_));
  NAND2_X1  g0583(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g0584(.A1(new_n784_), .A2(new_n424_), .A3(new_n432_), .A4(new_n779_), .ZN(new_n785_));
  NAND2_X1  g0585(.A1(new_n781_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g0586(.A(KEYINPUT63), .ZN(new_n787_));
  XNOR2_X1  g0587(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  NAND2_X1  g0588(.A1(new_n683_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g0589(.A1(new_n694_), .A2(new_n655_), .ZN(new_n790_));
  INV_X1    g0590(.A(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g0591(.A(new_n786_), .B(KEYINPUT63), .ZN(new_n792_));
  NAND3_X1  g0592(.A1(new_n792_), .A2(new_n672_), .A3(new_n682_), .ZN(new_n793_));
  NAND3_X1  g0593(.A1(new_n789_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g0594(.A(KEYINPUT65), .ZN(new_n795_));
  NAND2_X1  g0595(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OR2_X1    g0596(.A1(new_n794_), .A2(new_n795_), .ZN(new_n797_));
  NAND2_X1  g0597(.A1(new_n789_), .A2(new_n793_), .ZN(new_n798_));
  NAND2_X1  g0598(.A1(new_n798_), .A2(new_n790_), .ZN(new_n799_));
  NAND2_X1  g0599(.A1(new_n799_), .A2(KEYINPUT64), .ZN(new_n800_));
  INV_X1    g0600(.A(KEYINPUT64), .ZN(new_n801_));
  NAND3_X1  g0601(.A1(new_n798_), .A2(new_n801_), .A3(new_n790_), .ZN(new_n802_));
  AOI22_X1  g0602(.A1(new_n796_), .A2(new_n797_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g0603(.A(new_n704_), .ZN(new_n804_));
  OAI21_X1  g0604(.A(KEYINPUT66), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g0605(.A1(new_n797_), .A2(new_n796_), .ZN(new_n806_));
  NAND2_X1  g0606(.A1(new_n800_), .A2(new_n802_), .ZN(new_n807_));
  NAND2_X1  g0607(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g0608(.A(KEYINPUT66), .ZN(new_n809_));
  NAND3_X1  g0609(.A1(new_n808_), .A2(new_n809_), .A3(new_n704_), .ZN(new_n810_));
  NAND2_X1  g0610(.A1(new_n805_), .A2(new_n810_), .ZN(new_n811_));
  AOI22_X1  g0611(.A1(G137), .A2(new_n717_), .B1(new_n718_), .B2(G143), .ZN(new_n812_));
  INV_X1    g0612(.A(G150), .ZN(new_n813_));
  INV_X1    g0613(.A(G159), .ZN(new_n814_));
  OAI221_X1 g0614(.A(new_n812_), .B1(new_n813_), .B2(new_n724_), .C1(new_n814_), .C2(new_n725_), .ZN(new_n815_));
  XNOR2_X1  g0615(.A(new_n815_), .B(KEYINPUT68), .ZN(new_n816_));
  AOI21_X1  g0616(.A(KEYINPUT67), .B1(new_n747_), .B2(G50), .ZN(new_n817_));
  AND3_X1   g0617(.A1(new_n747_), .A2(KEYINPUT67), .A3(G50), .ZN(new_n818_));
  OAI221_X1 g0618(.A(new_n816_), .B1(new_n223_), .B2(new_n738_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g0619(.A(new_n819_), .B(KEYINPUT69), .ZN(new_n820_));
  NOR2_X1   g0620(.A1(new_n743_), .A2(new_n213_), .ZN(new_n821_));
  AOI211_X1 g0621(.A(G33), .B(new_n821_), .C1(new_n740_), .C2(G132), .ZN(new_n822_));
  NAND2_X1  g0622(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g0623(.A(G294), .ZN(new_n824_));
  OAI22_X1  g0624(.A1(new_n745_), .A2(new_n824_), .B1(new_n569_), .B2(new_n724_), .ZN(new_n825_));
  AOI211_X1 g0625(.A(new_n825_), .B(new_n739_), .C1(G303), .C2(new_n717_), .ZN(new_n826_));
  NAND2_X1  g0626(.A1(new_n728_), .A2(G87), .ZN(new_n827_));
  OAI21_X1  g0627(.A(G33), .B1(new_n725_), .B2(new_n579_), .ZN(new_n828_));
  AOI21_X1  g0628(.A(new_n828_), .B1(G107), .B2(new_n747_), .ZN(new_n829_));
  NAND2_X1  g0629(.A1(new_n740_), .A2(G311), .ZN(new_n830_));
  NAND4_X1  g0630(.A1(new_n826_), .A2(new_n827_), .A3(new_n829_), .A4(new_n830_), .ZN(new_n831_));
  AOI21_X1  g0631(.A(new_n710_), .B1(new_n823_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g0632(.A1(new_n709_), .A2(new_n761_), .ZN(new_n833_));
  AOI211_X1 g0633(.A(new_n775_), .B(new_n832_), .C1(new_n202_), .C2(new_n833_), .ZN(new_n834_));
  OR2_X1    g0634(.A1(new_n786_), .A2(new_n762_), .ZN(new_n835_));
  NAND2_X1  g0635(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g0636(.A(new_n665_), .ZN(new_n837_));
  OAI21_X1  g0637(.A(new_n836_), .B1(new_n803_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g0638(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g0639(.A1(new_n811_), .A2(new_n839_), .ZN(G384));
  OAI21_X1  g0640(.A(new_n500_), .B1(new_n229_), .B2(new_n219_), .ZN(new_n841_));
  NOR2_X1   g0641(.A1(new_n211_), .A2(new_n579_), .ZN(new_n842_));
  OAI21_X1  g0642(.A(G77), .B1(new_n223_), .B2(new_n213_), .ZN(new_n843_));
  OAI22_X1  g0643(.A1(new_n843_), .A2(new_n208_), .B1(G50), .B2(new_n213_), .ZN(new_n844_));
  NOR2_X1   g0644(.A1(new_n264_), .A2(G13), .ZN(new_n845_));
  AOI22_X1  g0645(.A1(new_n841_), .A2(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g0646(.A(new_n638_), .B(KEYINPUT70), .ZN(new_n847_));
  INV_X1    g0647(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g0648(.A1(new_n305_), .A2(KEYINPUT71), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g0649(.A(KEYINPUT71), .ZN(new_n850_));
  OAI21_X1  g0650(.A(new_n850_), .B1(new_n311_), .B2(new_n847_), .ZN(new_n851_));
  NAND2_X1  g0651(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g0652(.A(new_n852_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n853_));
  NAND3_X1  g0653(.A1(new_n274_), .A2(new_n269_), .A3(new_n847_), .ZN(new_n854_));
  NAND2_X1  g0654(.A1(new_n305_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g0655(.A(new_n310_), .ZN(new_n856_));
  NAND2_X1  g0656(.A1(new_n305_), .A2(KEYINPUT72), .ZN(new_n857_));
  INV_X1    g0657(.A(KEYINPUT72), .ZN(new_n858_));
  NAND2_X1  g0658(.A1(new_n311_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g0659(.A(new_n856_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g0660(.A(KEYINPUT73), .ZN(new_n861_));
  OAI21_X1  g0661(.A(new_n855_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  AOI211_X1 g0662(.A(KEYINPUT73), .B(new_n856_), .C1(new_n857_), .C2(new_n859_), .ZN(new_n863_));
  OAI21_X1  g0663(.A(new_n853_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g0664(.A1(new_n378_), .A2(new_n642_), .ZN(new_n865_));
  NAND3_X1  g0665(.A1(new_n377_), .A2(new_n382_), .A3(new_n865_), .ZN(new_n866_));
  OAI211_X1 g0666(.A(new_n380_), .B(new_n375_), .C1(new_n378_), .C2(new_n642_), .ZN(new_n867_));
  NAND2_X1  g0667(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g0668(.A1(new_n864_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g0669(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g0670(.A1(new_n870_), .A2(new_n786_), .ZN(new_n871_));
  NAND3_X1  g0671(.A1(new_n437_), .A2(new_n695_), .A3(new_n871_), .ZN(new_n872_));
  NOR2_X1   g0672(.A1(new_n871_), .A2(new_n694_), .ZN(new_n873_));
  INV_X1    g0673(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g0674(.A(new_n872_), .B1(new_n874_), .B2(new_n437_), .ZN(new_n875_));
  INV_X1    g0675(.A(KEYINPUT75), .ZN(new_n876_));
  NAND2_X1  g0676(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g0677(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g0678(.A1(new_n875_), .A2(new_n876_), .ZN(new_n879_));
  NOR3_X1   g0679(.A1(new_n878_), .A2(new_n655_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g0680(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g0681(.A1(new_n375_), .A2(new_n641_), .ZN(new_n882_));
  NAND2_X1  g0682(.A1(new_n864_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g0683(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g0684(.A1(new_n306_), .A2(new_n848_), .ZN(new_n885_));
  INV_X1    g0685(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g0686(.A1(new_n429_), .A2(new_n641_), .ZN(new_n887_));
  AOI21_X1  g0687(.A(new_n641_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n888_));
  AOI21_X1  g0688(.A(new_n887_), .B1(new_n888_), .B2(new_n786_), .ZN(new_n889_));
  OAI211_X1 g0689(.A(KEYINPUT74), .B(new_n886_), .C1(new_n889_), .C2(new_n869_), .ZN(new_n890_));
  INV_X1    g0690(.A(KEYINPUT74), .ZN(new_n891_));
  OAI211_X1 g0691(.A(new_n786_), .B(new_n642_), .C1(new_n674_), .C2(new_n680_), .ZN(new_n892_));
  INV_X1    g0692(.A(new_n887_), .ZN(new_n893_));
  AOI21_X1  g0693(.A(new_n869_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g0694(.A(new_n891_), .B1(new_n894_), .B2(new_n885_), .ZN(new_n895_));
  AOI21_X1  g0695(.A(new_n884_), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g0696(.A1(new_n437_), .A2(new_n683_), .ZN(new_n897_));
  NAND2_X1  g0697(.A1(new_n897_), .A2(new_n619_), .ZN(new_n898_));
  XOR2_X1   g0698(.A(new_n896_), .B(new_n898_), .Z(new_n899_));
  OAI22_X1  g0699(.A1(new_n881_), .A2(new_n899_), .B1(new_n264_), .B2(new_n702_), .ZN(new_n900_));
  INV_X1    g0700(.A(new_n899_), .ZN(new_n901_));
  NOR2_X1   g0701(.A1(new_n901_), .A2(new_n880_), .ZN(new_n902_));
  OAI21_X1  g0702(.A(new_n846_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  XOR2_X1   g0703(.A(new_n903_), .B(KEYINPUT76), .Z(G367));
  NAND2_X1  g0704(.A1(new_n520_), .A2(new_n641_), .ZN(new_n905_));
  OR2_X1    g0705(.A1(new_n472_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g0706(.A1(new_n472_), .A2(new_n524_), .A3(new_n905_), .ZN(new_n907_));
  NAND2_X1  g0707(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g0708(.A(new_n908_), .ZN(new_n909_));
  INV_X1    g0709(.A(new_n621_), .ZN(new_n910_));
  NAND2_X1  g0710(.A1(new_n513_), .A2(new_n641_), .ZN(new_n911_));
  XOR2_X1   g0711(.A(new_n517_), .B(new_n911_), .Z(new_n912_));
  OAI21_X1  g0712(.A(new_n910_), .B1(new_n659_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g0713(.A(new_n909_), .B1(new_n913_), .B2(new_n642_), .ZN(new_n914_));
  XNOR2_X1  g0714(.A(new_n914_), .B(KEYINPUT79), .ZN(new_n915_));
  INV_X1    g0715(.A(new_n915_), .ZN(new_n916_));
  NAND3_X1  g0716(.A1(new_n913_), .A2(new_n642_), .A3(new_n909_), .ZN(new_n917_));
  OR2_X1    g0717(.A1(new_n917_), .A2(KEYINPUT77), .ZN(new_n918_));
  NAND2_X1  g0718(.A1(new_n917_), .A2(KEYINPUT77), .ZN(new_n919_));
  NAND3_X1  g0719(.A1(new_n644_), .A2(G330), .A3(new_n654_), .ZN(new_n920_));
  NOR2_X1   g0720(.A1(new_n920_), .A2(new_n912_), .ZN(new_n921_));
  XNOR2_X1  g0721(.A(new_n921_), .B(KEYINPUT78), .ZN(new_n922_));
  AOI22_X1  g0722(.A1(new_n918_), .A2(new_n919_), .B1(new_n922_), .B2(KEYINPUT80), .ZN(new_n923_));
  OAI211_X1 g0723(.A(new_n916_), .B(new_n923_), .C1(KEYINPUT80), .C2(new_n922_), .ZN(new_n924_));
  INV_X1    g0724(.A(KEYINPUT80), .ZN(new_n925_));
  INV_X1    g0725(.A(new_n922_), .ZN(new_n926_));
  AND2_X1   g0726(.A1(new_n918_), .A2(new_n919_), .ZN(new_n927_));
  OAI211_X1 g0727(.A(new_n925_), .B(new_n926_), .C1(new_n927_), .C2(new_n915_), .ZN(new_n928_));
  AND2_X1   g0728(.A1(new_n924_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g0729(.A1(new_n644_), .A2(G330), .ZN(new_n930_));
  NAND3_X1  g0730(.A1(new_n930_), .A2(new_n653_), .A3(new_n652_), .ZN(new_n931_));
  NAND2_X1  g0731(.A1(new_n931_), .A2(new_n920_), .ZN(new_n932_));
  NOR2_X1   g0732(.A1(new_n634_), .A2(new_n641_), .ZN(new_n933_));
  XOR2_X1   g0733(.A(new_n932_), .B(new_n933_), .Z(new_n934_));
  INV_X1    g0734(.A(new_n934_), .ZN(new_n935_));
  NAND2_X1  g0735(.A1(new_n935_), .A2(new_n696_), .ZN(new_n936_));
  INV_X1    g0736(.A(KEYINPUT84), .ZN(new_n937_));
  INV_X1    g0737(.A(new_n912_), .ZN(new_n938_));
  OAI21_X1  g0738(.A(new_n938_), .B1(new_n659_), .B2(new_n641_), .ZN(new_n939_));
  INV_X1    g0739(.A(KEYINPUT83), .ZN(new_n940_));
  XNOR2_X1  g0740(.A(new_n939_), .B(new_n940_), .ZN(new_n941_));
  INV_X1    g0741(.A(new_n517_), .ZN(new_n942_));
  OAI211_X1 g0742(.A(new_n942_), .B(new_n642_), .C1(new_n658_), .C2(new_n625_), .ZN(new_n943_));
  XOR2_X1   g0743(.A(new_n943_), .B(KEYINPUT82), .Z(new_n944_));
  XOR2_X1   g0744(.A(new_n657_), .B(KEYINPUT81), .Z(new_n945_));
  NAND3_X1  g0745(.A1(new_n941_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  INV_X1    g0746(.A(new_n946_), .ZN(new_n947_));
  AOI21_X1  g0747(.A(new_n945_), .B1(new_n941_), .B2(new_n944_), .ZN(new_n948_));
  OAI21_X1  g0748(.A(new_n937_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  INV_X1    g0749(.A(new_n948_), .ZN(new_n950_));
  NAND3_X1  g0750(.A1(new_n950_), .A2(KEYINPUT84), .A3(new_n946_), .ZN(new_n951_));
  AOI21_X1  g0751(.A(new_n936_), .B1(new_n949_), .B2(new_n951_), .ZN(new_n952_));
  XOR2_X1   g0752(.A(new_n696_), .B(KEYINPUT85), .Z(new_n953_));
  OAI211_X1 g0753(.A(new_n929_), .B(new_n665_), .C1(new_n952_), .C2(new_n953_), .ZN(new_n954_));
  NAND3_X1  g0754(.A1(new_n924_), .A2(new_n928_), .A3(new_n704_), .ZN(new_n955_));
  INV_X1    g0755(.A(KEYINPUT87), .ZN(new_n956_));
  AOI21_X1  g0756(.A(new_n253_), .B1(new_n756_), .B2(G283), .ZN(new_n957_));
  NAND2_X1  g0757(.A1(new_n728_), .A2(G97), .ZN(new_n958_));
  OAI211_X1 g0758(.A(new_n957_), .B(new_n958_), .C1(new_n579_), .C2(new_n731_), .ZN(new_n959_));
  INV_X1    g0759(.A(new_n724_), .ZN(new_n960_));
  AOI22_X1  g0760(.A1(new_n960_), .A2(G294), .B1(G311), .B2(new_n717_), .ZN(new_n961_));
  OAI221_X1 g0761(.A(new_n961_), .B1(new_n219_), .B2(new_n738_), .C1(new_n585_), .C2(new_n745_), .ZN(new_n962_));
  AOI211_X1 g0762(.A(new_n959_), .B(new_n962_), .C1(G317), .C2(new_n740_), .ZN(new_n963_));
  AOI21_X1  g0763(.A(G33), .B1(new_n960_), .B2(G159), .ZN(new_n964_));
  OAI221_X1 g0764(.A(new_n964_), .B1(new_n223_), .B2(new_n731_), .C1(new_n202_), .C2(new_n743_), .ZN(new_n965_));
  AOI22_X1  g0765(.A1(new_n756_), .A2(G50), .B1(G150), .B2(new_n718_), .ZN(new_n966_));
  INV_X1    g0766(.A(G143), .ZN(new_n967_));
  OAI221_X1 g0767(.A(new_n966_), .B1(new_n213_), .B2(new_n738_), .C1(new_n967_), .C2(new_n752_), .ZN(new_n968_));
  AOI211_X1 g0768(.A(new_n965_), .B(new_n968_), .C1(G137), .C2(new_n740_), .ZN(new_n969_));
  OAI21_X1  g0769(.A(new_n709_), .B1(new_n963_), .B2(new_n969_), .ZN(new_n970_));
  NAND2_X1  g0770(.A1(new_n238_), .A2(new_n766_), .ZN(new_n971_));
  AOI21_X1  g0771(.A(new_n765_), .B1(new_n662_), .B2(new_n387_), .ZN(new_n972_));
  AOI21_X1  g0772(.A(new_n775_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  OAI211_X1 g0773(.A(new_n970_), .B(new_n973_), .C1(new_n908_), .C2(new_n764_), .ZN(new_n974_));
  XOR2_X1   g0774(.A(new_n974_), .B(KEYINPUT86), .Z(new_n975_));
  AND3_X1   g0775(.A1(new_n955_), .A2(new_n956_), .A3(new_n975_), .ZN(new_n976_));
  AOI21_X1  g0776(.A(new_n956_), .B1(new_n955_), .B2(new_n975_), .ZN(new_n977_));
  OAI21_X1  g0777(.A(new_n954_), .B1(new_n976_), .B2(new_n977_), .ZN(new_n978_));
  XNOR2_X1  g0778(.A(new_n978_), .B(KEYINPUT88), .ZN(G387));
  NAND2_X1  g0779(.A1(new_n953_), .A2(new_n934_), .ZN(new_n980_));
  XNOR2_X1  g0780(.A(new_n980_), .B(KEYINPUT89), .ZN(new_n981_));
  NAND3_X1  g0781(.A1(new_n981_), .A2(new_n665_), .A3(new_n936_), .ZN(new_n982_));
  INV_X1    g0782(.A(new_n771_), .ZN(new_n983_));
  NOR2_X1   g0783(.A1(new_n442_), .A2(G116), .ZN(new_n984_));
  OAI22_X1  g0784(.A1(new_n983_), .A2(new_n984_), .B1(G107), .B2(new_n206_), .ZN(new_n985_));
  OAI21_X1  g0785(.A(new_n451_), .B1(new_n213_), .B2(new_n202_), .ZN(new_n986_));
  NOR3_X1   g0786(.A1(new_n986_), .A2(G50), .A3(new_n223_), .ZN(new_n987_));
  AOI21_X1  g0787(.A(new_n767_), .B1(new_n987_), .B2(new_n984_), .ZN(new_n988_));
  NAND2_X1  g0788(.A1(new_n241_), .A2(G45), .ZN(new_n989_));
  AOI21_X1  g0789(.A(new_n985_), .B1(new_n988_), .B2(new_n989_), .ZN(new_n990_));
  OAI21_X1  g0790(.A(new_n774_), .B1(new_n990_), .B2(new_n765_), .ZN(new_n991_));
  AOI22_X1  g0791(.A1(G159), .A2(new_n717_), .B1(new_n718_), .B2(G50), .ZN(new_n992_));
  OAI21_X1  g0792(.A(new_n992_), .B1(new_n213_), .B2(new_n725_), .ZN(new_n993_));
  AOI21_X1  g0793(.A(G33), .B1(new_n960_), .B2(G58), .ZN(new_n994_));
  OAI211_X1 g0794(.A(new_n994_), .B(new_n958_), .C1(new_n202_), .C2(new_n731_), .ZN(new_n995_));
  AOI211_X1 g0795(.A(new_n993_), .B(new_n995_), .C1(G150), .C2(new_n740_), .ZN(new_n996_));
  NAND2_X1  g0796(.A1(new_n737_), .A2(new_n387_), .ZN(new_n997_));
  XNOR2_X1  g0797(.A(new_n997_), .B(KEYINPUT90), .ZN(new_n998_));
  AOI22_X1  g0798(.A1(G322), .A2(new_n717_), .B1(new_n718_), .B2(G317), .ZN(new_n999_));
  XNOR2_X1  g0799(.A(new_n999_), .B(KEYINPUT91), .ZN(new_n1000_));
  NAND2_X1  g0800(.A1(new_n960_), .A2(new_n757_), .ZN(new_n1001_));
  OAI211_X1 g0801(.A(new_n1001_), .B(G33), .C1(new_n585_), .C2(new_n725_), .ZN(new_n1002_));
  INV_X1    g0802(.A(new_n740_), .ZN(new_n1003_));
  OAI22_X1  g0803(.A1(new_n569_), .A2(new_n738_), .B1(new_n1003_), .B2(new_n753_), .ZN(new_n1004_));
  OAI22_X1  g0804(.A1(new_n743_), .A2(new_n579_), .B1(new_n731_), .B2(new_n824_), .ZN(new_n1005_));
  NOR3_X1   g0805(.A1(new_n1002_), .A2(new_n1004_), .A3(new_n1005_), .ZN(new_n1006_));
  AOI22_X1  g0806(.A1(new_n996_), .A2(new_n998_), .B1(new_n1000_), .B2(new_n1006_), .ZN(new_n1007_));
  OR2_X1    g0807(.A1(new_n1007_), .A2(KEYINPUT92), .ZN(new_n1008_));
  AOI21_X1  g0808(.A(new_n710_), .B1(new_n1007_), .B2(KEYINPUT92), .ZN(new_n1009_));
  AOI21_X1  g0809(.A(new_n991_), .B1(new_n1008_), .B2(new_n1009_), .ZN(new_n1010_));
  OAI21_X1  g0810(.A(new_n1010_), .B1(new_n654_), .B2(new_n764_), .ZN(new_n1011_));
  OAI21_X1  g0811(.A(new_n1011_), .B1(new_n934_), .B2(new_n703_), .ZN(new_n1012_));
  INV_X1    g0812(.A(new_n1012_), .ZN(new_n1013_));
  NAND2_X1  g0813(.A1(new_n982_), .A2(new_n1013_), .ZN(G393));
  AND3_X1   g0814(.A1(new_n936_), .A2(new_n946_), .A3(new_n950_), .ZN(new_n1015_));
  NOR3_X1   g0815(.A1(new_n952_), .A2(new_n837_), .A3(new_n1015_), .ZN(new_n1016_));
  NAND2_X1  g0816(.A1(new_n949_), .A2(new_n951_), .ZN(new_n1017_));
  NAND2_X1  g0817(.A1(new_n1017_), .A2(new_n704_), .ZN(new_n1018_));
  AOI21_X1  g0818(.A(new_n765_), .B1(new_n229_), .B2(new_n662_), .ZN(new_n1019_));
  NAND2_X1  g0819(.A1(new_n245_), .A2(new_n766_), .ZN(new_n1020_));
  AOI21_X1  g0820(.A(new_n775_), .B1(new_n1019_), .B2(new_n1020_), .ZN(new_n1021_));
  NAND2_X1  g0821(.A1(new_n737_), .A2(G77), .ZN(new_n1022_));
  XOR2_X1   g0822(.A(new_n1022_), .B(KEYINPUT93), .Z(new_n1023_));
  AOI21_X1  g0823(.A(G33), .B1(new_n960_), .B2(G50), .ZN(new_n1024_));
  OAI211_X1 g0824(.A(new_n1024_), .B(new_n827_), .C1(new_n213_), .C2(new_n731_), .ZN(new_n1025_));
  AOI22_X1  g0825(.A1(G150), .A2(new_n717_), .B1(new_n718_), .B2(G159), .ZN(new_n1026_));
  OAI221_X1 g0826(.A(new_n1026_), .B1(new_n223_), .B2(new_n725_), .C1(new_n967_), .C2(new_n1003_), .ZN(new_n1027_));
  OR3_X1    g0827(.A1(new_n1023_), .A2(new_n1025_), .A3(new_n1027_), .ZN(new_n1028_));
  AND2_X1   g0828(.A1(new_n1028_), .A2(KEYINPUT94), .ZN(new_n1029_));
  NOR2_X1   g0829(.A1(new_n1028_), .A2(KEYINPUT94), .ZN(new_n1030_));
  AOI21_X1  g0830(.A(new_n253_), .B1(new_n756_), .B2(G294), .ZN(new_n1031_));
  OAI211_X1 g0831(.A(new_n1031_), .B(new_n729_), .C1(new_n569_), .C2(new_n731_), .ZN(new_n1032_));
  AOI22_X1  g0832(.A1(new_n960_), .A2(G303), .B1(G311), .B2(new_n718_), .ZN(new_n1033_));
  OAI221_X1 g0833(.A(new_n1033_), .B1(new_n754_), .B2(new_n752_), .C1(new_n744_), .C2(new_n1003_), .ZN(new_n1034_));
  AOI211_X1 g0834(.A(new_n1032_), .B(new_n1034_), .C1(G116), .C2(new_n737_), .ZN(new_n1035_));
  NOR3_X1   g0835(.A1(new_n1029_), .A2(new_n1030_), .A3(new_n1035_), .ZN(new_n1036_));
  OAI221_X1 g0836(.A(new_n1021_), .B1(new_n1036_), .B2(new_n710_), .C1(new_n938_), .C2(new_n764_), .ZN(new_n1037_));
  NAND2_X1  g0837(.A1(new_n1018_), .A2(new_n1037_), .ZN(new_n1038_));
  OR2_X1    g0838(.A1(new_n1016_), .A2(new_n1038_), .ZN(G390));
  NAND4_X1  g0839(.A1(new_n692_), .A2(G330), .A3(new_n693_), .A4(new_n786_), .ZN(new_n1040_));
  INV_X1    g0840(.A(new_n868_), .ZN(new_n1041_));
  NOR2_X1   g0841(.A1(new_n1040_), .A2(new_n1041_), .ZN(new_n1042_));
  INV_X1    g0842(.A(new_n1042_), .ZN(new_n1043_));
  NAND2_X1  g0843(.A1(new_n887_), .A2(new_n868_), .ZN(new_n1044_));
  NAND2_X1  g0844(.A1(new_n1044_), .A2(KEYINPUT95), .ZN(new_n1045_));
  INV_X1    g0845(.A(KEYINPUT95), .ZN(new_n1046_));
  NAND3_X1  g0846(.A1(new_n887_), .A2(new_n868_), .A3(new_n1046_), .ZN(new_n1047_));
  AOI21_X1  g0847(.A(new_n882_), .B1(new_n1045_), .B2(new_n1047_), .ZN(new_n1048_));
  NAND4_X1  g0848(.A1(new_n630_), .A2(new_n642_), .A3(new_n786_), .A4(new_n868_), .ZN(new_n1049_));
  AND3_X1   g0849(.A1(new_n1048_), .A2(new_n864_), .A3(new_n1049_), .ZN(new_n1050_));
  AOI21_X1  g0850(.A(new_n864_), .B1(new_n1048_), .B2(new_n1049_), .ZN(new_n1051_));
  OAI21_X1  g0851(.A(new_n1043_), .B1(new_n1050_), .B2(new_n1051_), .ZN(new_n1052_));
  NAND2_X1  g0852(.A1(new_n1048_), .A2(new_n1049_), .ZN(new_n1053_));
  INV_X1    g0853(.A(new_n864_), .ZN(new_n1054_));
  NAND2_X1  g0854(.A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_));
  NAND3_X1  g0855(.A1(new_n1048_), .A2(new_n864_), .A3(new_n1049_), .ZN(new_n1056_));
  NAND3_X1  g0856(.A1(new_n1055_), .A2(new_n1056_), .A3(new_n1042_), .ZN(new_n1057_));
  AND2_X1   g0857(.A1(new_n1052_), .A2(new_n1057_), .ZN(new_n1058_));
  NAND3_X1  g0858(.A1(new_n695_), .A2(new_n656_), .A3(new_n788_), .ZN(new_n1059_));
  NAND2_X1  g0859(.A1(new_n892_), .A2(new_n893_), .ZN(new_n1060_));
  NAND2_X1  g0860(.A1(new_n1041_), .A2(KEYINPUT96), .ZN(new_n1061_));
  INV_X1    g0861(.A(new_n1061_), .ZN(new_n1062_));
  NOR2_X1   g0862(.A1(new_n1060_), .A2(new_n1062_), .ZN(new_n1063_));
  AOI21_X1  g0863(.A(new_n1061_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n1064_));
  NOR3_X1   g0864(.A1(new_n1059_), .A2(new_n1063_), .A3(new_n1064_), .ZN(new_n1065_));
  INV_X1    g0865(.A(new_n1065_), .ZN(new_n1066_));
  INV_X1    g0866(.A(KEYINPUT98), .ZN(new_n1067_));
  AND2_X1   g0867(.A1(new_n1040_), .A2(KEYINPUT97), .ZN(new_n1068_));
  NAND3_X1  g0868(.A1(new_n892_), .A2(new_n1041_), .A3(new_n893_), .ZN(new_n1069_));
  NAND3_X1  g0869(.A1(new_n1069_), .A2(new_n1049_), .A3(new_n1044_), .ZN(new_n1070_));
  NOR2_X1   g0870(.A1(new_n1068_), .A2(new_n1070_), .ZN(new_n1071_));
  NOR2_X1   g0871(.A1(new_n1040_), .A2(KEYINPUT97), .ZN(new_n1072_));
  INV_X1    g0872(.A(new_n1072_), .ZN(new_n1073_));
  AOI21_X1  g0873(.A(new_n1067_), .B1(new_n1071_), .B2(new_n1073_), .ZN(new_n1074_));
  INV_X1    g0874(.A(new_n892_), .ZN(new_n1075_));
  OAI21_X1  g0875(.A(new_n868_), .B1(new_n1075_), .B2(new_n887_), .ZN(new_n1076_));
  NAND2_X1  g0876(.A1(new_n1040_), .A2(KEYINPUT97), .ZN(new_n1077_));
  NAND3_X1  g0877(.A1(new_n1076_), .A2(new_n1077_), .A3(new_n1069_), .ZN(new_n1078_));
  NOR3_X1   g0878(.A1(new_n1078_), .A2(KEYINPUT98), .A3(new_n1072_), .ZN(new_n1079_));
  OAI21_X1  g0879(.A(new_n1066_), .B1(new_n1074_), .B2(new_n1079_), .ZN(new_n1080_));
  NAND2_X1  g0880(.A1(new_n1080_), .A2(KEYINPUT99), .ZN(new_n1081_));
  OAI21_X1  g0881(.A(KEYINPUT98), .B1(new_n1078_), .B2(new_n1072_), .ZN(new_n1082_));
  INV_X1    g0882(.A(new_n1070_), .ZN(new_n1083_));
  NAND4_X1  g0883(.A1(new_n1083_), .A2(new_n1073_), .A3(new_n1067_), .A4(new_n1077_), .ZN(new_n1084_));
  NAND2_X1  g0884(.A1(new_n1082_), .A2(new_n1084_), .ZN(new_n1085_));
  INV_X1    g0885(.A(KEYINPUT99), .ZN(new_n1086_));
  NAND3_X1  g0886(.A1(new_n1085_), .A2(new_n1086_), .A3(new_n1066_), .ZN(new_n1087_));
  NAND2_X1  g0887(.A1(new_n1081_), .A2(new_n1087_), .ZN(new_n1088_));
  NAND3_X1  g0888(.A1(new_n437_), .A2(new_n656_), .A3(new_n695_), .ZN(new_n1089_));
  NAND3_X1  g0889(.A1(new_n1089_), .A2(new_n619_), .A3(new_n897_), .ZN(new_n1090_));
  INV_X1    g0890(.A(KEYINPUT100), .ZN(new_n1091_));
  NAND2_X1  g0891(.A1(new_n1090_), .A2(new_n1091_), .ZN(new_n1092_));
  NAND4_X1  g0892(.A1(new_n1089_), .A2(new_n897_), .A3(new_n619_), .A4(KEYINPUT100), .ZN(new_n1093_));
  NAND2_X1  g0893(.A1(new_n1092_), .A2(new_n1093_), .ZN(new_n1094_));
  INV_X1    g0894(.A(new_n1094_), .ZN(new_n1095_));
  AOI21_X1  g0895(.A(new_n1058_), .B1(new_n1088_), .B2(new_n1095_), .ZN(new_n1096_));
  AOI21_X1  g0896(.A(new_n1086_), .B1(new_n1085_), .B2(new_n1066_), .ZN(new_n1097_));
  AOI211_X1 g0897(.A(KEYINPUT99), .B(new_n1065_), .C1(new_n1082_), .C2(new_n1084_), .ZN(new_n1098_));
  OAI211_X1 g0898(.A(new_n1058_), .B(new_n1095_), .C1(new_n1097_), .C2(new_n1098_), .ZN(new_n1099_));
  INV_X1    g0899(.A(new_n1099_), .ZN(new_n1100_));
  OAI21_X1  g0900(.A(new_n665_), .B1(new_n1096_), .B2(new_n1100_), .ZN(new_n1101_));
  NAND2_X1  g0901(.A1(new_n1052_), .A2(new_n1057_), .ZN(new_n1102_));
  NAND2_X1  g0902(.A1(new_n1102_), .A2(new_n704_), .ZN(new_n1103_));
  INV_X1    g0903(.A(KEYINPUT105), .ZN(new_n1104_));
  NAND2_X1  g0904(.A1(new_n1054_), .A2(new_n761_), .ZN(new_n1105_));
  XOR2_X1   g0905(.A(new_n1105_), .B(KEYINPUT104), .Z(new_n1106_));
  AOI21_X1  g0906(.A(new_n775_), .B1(new_n223_), .B2(new_n833_), .ZN(new_n1107_));
  AOI22_X1  g0907(.A1(G137), .A2(new_n960_), .B1(new_n756_), .B2(G143), .ZN(new_n1108_));
  INV_X1    g0908(.A(G132), .ZN(new_n1109_));
  OAI221_X1 g0909(.A(new_n1108_), .B1(new_n1109_), .B2(new_n745_), .C1(new_n814_), .C2(new_n738_), .ZN(new_n1110_));
  NAND2_X1  g0910(.A1(new_n740_), .A2(G125), .ZN(new_n1111_));
  XNOR2_X1  g0911(.A(new_n1111_), .B(KEYINPUT101), .ZN(new_n1112_));
  AOI21_X1  g0912(.A(G33), .B1(new_n717_), .B2(G128), .ZN(new_n1113_));
  OAI221_X1 g0913(.A(new_n1113_), .B1(new_n813_), .B2(new_n731_), .C1(new_n227_), .C2(new_n743_), .ZN(new_n1114_));
  NOR3_X1   g0914(.A1(new_n1110_), .A2(new_n1112_), .A3(new_n1114_), .ZN(new_n1115_));
  AOI22_X1  g0915(.A1(G283), .A2(new_n717_), .B1(new_n718_), .B2(G116), .ZN(new_n1116_));
  NAND2_X1  g0916(.A1(new_n960_), .A2(new_n548_), .ZN(new_n1117_));
  OAI211_X1 g0917(.A(new_n1116_), .B(new_n1117_), .C1(new_n230_), .C2(new_n725_), .ZN(new_n1118_));
  NOR3_X1   g0918(.A1(new_n1023_), .A2(new_n732_), .A3(new_n1118_), .ZN(new_n1119_));
  XOR2_X1   g0919(.A(new_n1119_), .B(KEYINPUT102), .Z(new_n1120_));
  OR3_X1    g0920(.A1(new_n1003_), .A2(KEYINPUT103), .A3(new_n824_), .ZN(new_n1121_));
  OAI21_X1  g0921(.A(KEYINPUT103), .B1(new_n1003_), .B2(new_n824_), .ZN(new_n1122_));
  AOI211_X1 g0922(.A(new_n253_), .B(new_n821_), .C1(new_n1121_), .C2(new_n1122_), .ZN(new_n1123_));
  AOI21_X1  g0923(.A(new_n1115_), .B1(new_n1120_), .B2(new_n1123_), .ZN(new_n1124_));
  OAI21_X1  g0924(.A(new_n1107_), .B1(new_n1124_), .B2(new_n710_), .ZN(new_n1125_));
  NOR2_X1   g0925(.A1(new_n1106_), .A2(new_n1125_), .ZN(new_n1126_));
  INV_X1    g0926(.A(new_n1126_), .ZN(new_n1127_));
  NAND3_X1  g0927(.A1(new_n1103_), .A2(new_n1104_), .A3(new_n1127_), .ZN(new_n1128_));
  AOI21_X1  g0928(.A(new_n804_), .B1(new_n1052_), .B2(new_n1057_), .ZN(new_n1129_));
  OAI21_X1  g0929(.A(KEYINPUT105), .B1(new_n1129_), .B2(new_n1126_), .ZN(new_n1130_));
  NAND2_X1  g0930(.A1(new_n1128_), .A2(new_n1130_), .ZN(new_n1131_));
  NAND2_X1  g0931(.A1(new_n1101_), .A2(new_n1131_), .ZN(G378));
  AOI22_X1  g0932(.A1(new_n756_), .A2(G137), .B1(G125), .B2(new_n717_), .ZN(new_n1133_));
  OAI221_X1 g0933(.A(new_n1133_), .B1(new_n1109_), .B2(new_n724_), .C1(new_n813_), .C2(new_n738_), .ZN(new_n1134_));
  AOI21_X1  g0934(.A(new_n1134_), .B1(G124), .B2(new_n740_), .ZN(new_n1135_));
  AOI211_X1 g0935(.A(G33), .B(G41), .C1(new_n718_), .C2(G128), .ZN(new_n1136_));
  OAI21_X1  g0936(.A(new_n1136_), .B1(new_n967_), .B2(new_n731_), .ZN(new_n1137_));
  AOI21_X1  g0937(.A(new_n1137_), .B1(G159), .B2(new_n728_), .ZN(new_n1138_));
  NAND2_X1  g0938(.A1(new_n473_), .A2(G33), .ZN(new_n1139_));
  XNOR2_X1  g0939(.A(new_n1139_), .B(KEYINPUT112), .ZN(new_n1140_));
  AOI21_X1  g0940(.A(G50), .B1(new_n253_), .B2(new_n473_), .ZN(new_n1141_));
  AOI22_X1  g0941(.A1(new_n1135_), .A2(new_n1138_), .B1(new_n1140_), .B2(new_n1141_), .ZN(new_n1142_));
  AOI22_X1  g0942(.A1(G116), .A2(new_n717_), .B1(new_n718_), .B2(G107), .ZN(new_n1143_));
  OAI221_X1 g0943(.A(new_n1143_), .B1(new_n230_), .B2(new_n724_), .C1(new_n446_), .C2(new_n725_), .ZN(new_n1144_));
  XOR2_X1   g0944(.A(new_n1144_), .B(KEYINPUT111), .Z(new_n1145_));
  AOI22_X1  g0945(.A1(G68), .A2(new_n737_), .B1(new_n740_), .B2(G283), .ZN(new_n1146_));
  NOR2_X1   g0946(.A1(new_n743_), .A2(new_n223_), .ZN(new_n1147_));
  INV_X1    g0947(.A(new_n1147_), .ZN(new_n1148_));
  AOI21_X1  g0948(.A(new_n1140_), .B1(new_n747_), .B2(G77), .ZN(new_n1149_));
  NAND3_X1  g0949(.A1(new_n1146_), .A2(new_n1148_), .A3(new_n1149_), .ZN(new_n1150_));
  OAI21_X1  g0950(.A(new_n1142_), .B1(new_n1145_), .B2(new_n1150_), .ZN(new_n1151_));
  INV_X1    g0951(.A(new_n1151_), .ZN(new_n1152_));
  AOI21_X1  g0952(.A(new_n710_), .B1(new_n1152_), .B2(KEYINPUT113), .ZN(new_n1153_));
  OAI21_X1  g0953(.A(new_n1153_), .B1(KEYINPUT113), .B2(new_n1152_), .ZN(new_n1154_));
  AOI21_X1  g0954(.A(new_n775_), .B1(new_n227_), .B2(new_n833_), .ZN(new_n1155_));
  NAND2_X1  g0955(.A1(new_n343_), .A2(new_n848_), .ZN(new_n1156_));
  XNOR2_X1  g0956(.A(new_n345_), .B(new_n1156_), .ZN(new_n1157_));
  INV_X1    g0957(.A(new_n1157_), .ZN(new_n1158_));
  OAI211_X1 g0958(.A(new_n1154_), .B(new_n1155_), .C1(new_n1158_), .C2(new_n762_), .ZN(new_n1159_));
  NOR2_X1   g0959(.A1(new_n874_), .A2(new_n655_), .ZN(new_n1160_));
  XNOR2_X1  g0960(.A(new_n883_), .B(KEYINPUT106), .ZN(new_n1161_));
  NAND2_X1  g0961(.A1(new_n1060_), .A2(new_n870_), .ZN(new_n1162_));
  NAND4_X1  g0962(.A1(new_n1161_), .A2(new_n886_), .A3(new_n1162_), .A4(new_n1158_), .ZN(new_n1163_));
  OAI211_X1 g0963(.A(new_n1160_), .B(new_n1163_), .C1(new_n896_), .C2(new_n1158_), .ZN(new_n1164_));
  INV_X1    g0964(.A(new_n1164_), .ZN(new_n1165_));
  AOI21_X1  g0965(.A(KEYINPUT74), .B1(new_n1162_), .B2(new_n886_), .ZN(new_n1166_));
  NOR3_X1   g0966(.A1(new_n894_), .A2(new_n891_), .A3(new_n885_), .ZN(new_n1167_));
  OAI211_X1 g0967(.A(new_n883_), .B(new_n1158_), .C1(new_n1166_), .C2(new_n1167_), .ZN(new_n1168_));
  NAND2_X1  g0968(.A1(new_n1168_), .A2(KEYINPUT110), .ZN(new_n1169_));
  INV_X1    g0969(.A(KEYINPUT110), .ZN(new_n1170_));
  NAND3_X1  g0970(.A1(new_n896_), .A2(new_n1170_), .A3(new_n1158_), .ZN(new_n1171_));
  OAI21_X1  g0971(.A(new_n1161_), .B1(new_n1166_), .B2(new_n1167_), .ZN(new_n1172_));
  NAND2_X1  g0972(.A1(new_n1172_), .A2(new_n1157_), .ZN(new_n1173_));
  NAND3_X1  g0973(.A1(new_n1169_), .A2(new_n1171_), .A3(new_n1173_), .ZN(new_n1174_));
  XNOR2_X1  g0974(.A(new_n1160_), .B(KEYINPUT109), .ZN(new_n1175_));
  AOI21_X1  g0975(.A(new_n1165_), .B1(new_n1174_), .B2(new_n1175_), .ZN(new_n1176_));
  OAI21_X1  g0976(.A(new_n1159_), .B1(new_n1176_), .B2(new_n804_), .ZN(new_n1177_));
  NOR2_X1   g0977(.A1(new_n1058_), .A2(new_n1094_), .ZN(new_n1178_));
  OAI21_X1  g0978(.A(new_n1178_), .B1(new_n1097_), .B2(new_n1098_), .ZN(new_n1179_));
  NAND2_X1  g0979(.A1(new_n1179_), .A2(new_n1095_), .ZN(new_n1180_));
  OAI21_X1  g0980(.A(new_n1163_), .B1(new_n896_), .B2(new_n1158_), .ZN(new_n1181_));
  INV_X1    g0981(.A(new_n1160_), .ZN(new_n1182_));
  NAND2_X1  g0982(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1183_));
  NAND3_X1  g0983(.A1(new_n1183_), .A2(KEYINPUT107), .A3(new_n1164_), .ZN(new_n1184_));
  INV_X1    g0984(.A(KEYINPUT107), .ZN(new_n1185_));
  NAND3_X1  g0985(.A1(new_n1181_), .A2(new_n1185_), .A3(new_n1182_), .ZN(new_n1186_));
  AND2_X1   g0986(.A1(new_n1184_), .A2(new_n1186_), .ZN(new_n1187_));
  NAND3_X1  g0987(.A1(new_n1180_), .A2(new_n1187_), .A3(new_n665_), .ZN(new_n1188_));
  INV_X1    g0988(.A(KEYINPUT108), .ZN(new_n1189_));
  AOI21_X1  g0989(.A(new_n1177_), .B1(new_n1188_), .B2(new_n1189_), .ZN(new_n1190_));
  NAND4_X1  g0990(.A1(new_n1180_), .A2(new_n1187_), .A3(KEYINPUT108), .A4(new_n665_), .ZN(new_n1191_));
  AND2_X1   g0991(.A1(new_n1190_), .A2(new_n1191_), .ZN(new_n1192_));
  INV_X1    g0992(.A(new_n1192_), .ZN(G375));
  NAND3_X1  g0993(.A1(new_n1081_), .A2(new_n1087_), .A3(new_n1094_), .ZN(new_n1194_));
  OAI21_X1  g0994(.A(new_n1095_), .B1(new_n1097_), .B2(new_n1098_), .ZN(new_n1195_));
  NAND3_X1  g0995(.A1(new_n1194_), .A2(new_n1195_), .A3(new_n665_), .ZN(new_n1196_));
  XOR2_X1   g0996(.A(new_n1196_), .B(KEYINPUT114), .Z(new_n1197_));
  NAND2_X1  g0997(.A1(new_n1041_), .A2(new_n761_), .ZN(new_n1198_));
  NOR3_X1   g0998(.A1(new_n709_), .A2(G68), .A3(new_n761_), .ZN(new_n1199_));
  NOR2_X1   g0999(.A1(new_n1003_), .A2(new_n585_), .ZN(new_n1200_));
  OAI22_X1  g1000(.A1(new_n752_), .A2(new_n824_), .B1(new_n745_), .B2(new_n569_), .ZN(new_n1201_));
  AOI211_X1 g1001(.A(new_n1200_), .B(new_n1201_), .C1(new_n548_), .C2(new_n756_), .ZN(new_n1202_));
  OAI221_X1 g1002(.A(G33), .B1(new_n724_), .B2(new_n579_), .C1(new_n743_), .C2(new_n202_), .ZN(new_n1203_));
  AOI21_X1  g1003(.A(new_n1203_), .B1(G97), .B2(new_n747_), .ZN(new_n1204_));
  NAND3_X1  g1004(.A1(new_n1202_), .A2(new_n998_), .A3(new_n1204_), .ZN(new_n1205_));
  NOR2_X1   g1005(.A1(new_n731_), .A2(new_n814_), .ZN(new_n1206_));
  XNOR2_X1  g1006(.A(new_n1206_), .B(KEYINPUT115), .ZN(new_n1207_));
  AOI211_X1 g1007(.A(G33), .B(new_n1147_), .C1(G132), .C2(new_n717_), .ZN(new_n1208_));
  NAND2_X1  g1008(.A1(new_n756_), .A2(G150), .ZN(new_n1209_));
  AOI22_X1  g1009(.A1(new_n960_), .A2(G143), .B1(G137), .B2(new_n718_), .ZN(new_n1210_));
  AOI22_X1  g1010(.A1(G50), .A2(new_n737_), .B1(new_n740_), .B2(G128), .ZN(new_n1211_));
  NAND4_X1  g1011(.A1(new_n1208_), .A2(new_n1209_), .A3(new_n1210_), .A4(new_n1211_), .ZN(new_n1212_));
  OAI21_X1  g1012(.A(new_n1205_), .B1(new_n1207_), .B2(new_n1212_), .ZN(new_n1213_));
  AOI211_X1 g1013(.A(new_n775_), .B(new_n1199_), .C1(new_n1213_), .C2(new_n709_), .ZN(new_n1214_));
  AOI22_X1  g1014(.A1(new_n1088_), .A2(new_n704_), .B1(new_n1198_), .B2(new_n1214_), .ZN(new_n1215_));
  NAND2_X1  g1015(.A1(new_n1197_), .A2(new_n1215_), .ZN(G381));
  INV_X1    g1016(.A(G396), .ZN(new_n1217_));
  NAND3_X1  g1017(.A1(new_n982_), .A2(new_n1217_), .A3(new_n1013_), .ZN(new_n1218_));
  OR3_X1    g1018(.A1(G390), .A2(G384), .A3(new_n1218_), .ZN(new_n1219_));
  NOR4_X1   g1019(.A1(G387), .A2(new_n1219_), .A3(G378), .A4(G381), .ZN(new_n1220_));
  NAND2_X1  g1020(.A1(new_n1220_), .A2(new_n1192_), .ZN(G407));
  INV_X1    g1021(.A(G378), .ZN(new_n1222_));
  NAND3_X1  g1022(.A1(new_n1192_), .A2(new_n640_), .A3(new_n1222_), .ZN(new_n1223_));
  NAND3_X1  g1023(.A1(G407), .A2(G213), .A3(new_n1223_), .ZN(G409));
  NOR2_X1   g1024(.A1(new_n637_), .A2(G343), .ZN(new_n1225_));
  NOR2_X1   g1025(.A1(new_n1179_), .A2(new_n1176_), .ZN(new_n1226_));
  AND3_X1   g1026(.A1(new_n1184_), .A2(new_n1094_), .A3(new_n1186_), .ZN(new_n1227_));
  OAI21_X1  g1027(.A(new_n665_), .B1(new_n1226_), .B2(new_n1227_), .ZN(new_n1228_));
  INV_X1    g1028(.A(new_n1177_), .ZN(new_n1229_));
  AOI21_X1  g1029(.A(new_n1225_), .B1(new_n1228_), .B2(new_n1229_), .ZN(new_n1230_));
  INV_X1    g1030(.A(KEYINPUT117), .ZN(new_n1231_));
  NAND2_X1  g1031(.A1(new_n1195_), .A2(new_n1102_), .ZN(new_n1232_));
  AOI21_X1  g1032(.A(new_n837_), .B1(new_n1232_), .B2(new_n1099_), .ZN(new_n1233_));
  NAND2_X1  g1033(.A1(new_n1131_), .A2(KEYINPUT116), .ZN(new_n1234_));
  INV_X1    g1034(.A(KEYINPUT116), .ZN(new_n1235_));
  NAND3_X1  g1035(.A1(new_n1128_), .A2(new_n1235_), .A3(new_n1130_), .ZN(new_n1236_));
  NAND2_X1  g1036(.A1(new_n1234_), .A2(new_n1236_), .ZN(new_n1237_));
  OAI21_X1  g1037(.A(new_n1231_), .B1(new_n1233_), .B2(new_n1237_), .ZN(new_n1238_));
  INV_X1    g1038(.A(new_n1236_), .ZN(new_n1239_));
  AOI21_X1  g1039(.A(new_n1235_), .B1(new_n1128_), .B2(new_n1130_), .ZN(new_n1240_));
  NOR2_X1   g1040(.A1(new_n1239_), .A2(new_n1240_), .ZN(new_n1241_));
  NAND3_X1  g1041(.A1(new_n1101_), .A2(new_n1241_), .A3(KEYINPUT117), .ZN(new_n1242_));
  NAND3_X1  g1042(.A1(new_n1230_), .A2(new_n1238_), .A3(new_n1242_), .ZN(new_n1243_));
  INV_X1    g1043(.A(new_n1225_), .ZN(new_n1244_));
  NAND4_X1  g1044(.A1(new_n1190_), .A2(G378), .A3(new_n1191_), .A4(new_n1244_), .ZN(new_n1245_));
  AND2_X1   g1045(.A1(new_n1243_), .A2(new_n1245_), .ZN(new_n1246_));
  NAND2_X1  g1046(.A1(new_n1215_), .A2(new_n1196_), .ZN(new_n1247_));
  AOI21_X1  g1047(.A(new_n838_), .B1(new_n810_), .B2(new_n805_), .ZN(new_n1248_));
  NAND2_X1  g1048(.A1(new_n1247_), .A2(new_n1248_), .ZN(new_n1249_));
  NAND3_X1  g1049(.A1(G384), .A2(new_n1215_), .A3(new_n1196_), .ZN(new_n1250_));
  NAND2_X1  g1050(.A1(new_n1225_), .A2(G2897), .ZN(new_n1251_));
  INV_X1    g1051(.A(new_n1251_), .ZN(new_n1252_));
  AND3_X1   g1052(.A1(new_n1249_), .A2(new_n1250_), .A3(new_n1252_), .ZN(new_n1253_));
  NAND3_X1  g1053(.A1(new_n1246_), .A2(KEYINPUT125), .A3(new_n1253_), .ZN(new_n1254_));
  NAND2_X1  g1054(.A1(new_n1243_), .A2(new_n1245_), .ZN(new_n1255_));
  INV_X1    g1055(.A(KEYINPUT119), .ZN(new_n1256_));
  NAND2_X1  g1056(.A1(new_n1249_), .A2(new_n1250_), .ZN(new_n1257_));
  OAI21_X1  g1057(.A(new_n1256_), .B1(new_n1257_), .B2(new_n1252_), .ZN(new_n1258_));
  NAND4_X1  g1058(.A1(new_n1249_), .A2(new_n1250_), .A3(KEYINPUT119), .A4(new_n1251_), .ZN(new_n1259_));
  NAND3_X1  g1059(.A1(new_n1255_), .A2(new_n1258_), .A3(new_n1259_), .ZN(new_n1260_));
  NAND3_X1  g1060(.A1(new_n1243_), .A2(new_n1245_), .A3(new_n1253_), .ZN(new_n1261_));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262_));
  NAND2_X1  g1062(.A1(new_n1261_), .A2(new_n1262_), .ZN(new_n1263_));
  NAND3_X1  g1063(.A1(new_n1254_), .A2(new_n1260_), .A3(new_n1263_), .ZN(new_n1264_));
  NAND2_X1  g1064(.A1(new_n1264_), .A2(KEYINPUT126), .ZN(new_n1265_));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266_));
  NAND4_X1  g1066(.A1(new_n1254_), .A2(new_n1266_), .A3(new_n1260_), .A4(new_n1263_), .ZN(new_n1267_));
  AOI21_X1  g1067(.A(new_n1252_), .B1(new_n1249_), .B2(new_n1250_), .ZN(new_n1268_));
  AND3_X1   g1068(.A1(new_n1243_), .A2(new_n1245_), .A3(new_n1268_), .ZN(new_n1269_));
  AOI21_X1  g1069(.A(KEYINPUT118), .B1(new_n1257_), .B2(new_n1252_), .ZN(new_n1270_));
  INV_X1    g1070(.A(KEYINPUT118), .ZN(new_n1271_));
  AOI211_X1 g1071(.A(new_n1271_), .B(new_n1251_), .C1(new_n1249_), .C2(new_n1250_), .ZN(new_n1272_));
  NOR2_X1   g1072(.A1(new_n1270_), .A2(new_n1272_), .ZN(new_n1273_));
  AOI21_X1  g1073(.A(new_n1269_), .B1(new_n1255_), .B2(new_n1273_), .ZN(new_n1274_));
  NOR2_X1   g1074(.A1(new_n1016_), .A2(new_n1038_), .ZN(new_n1275_));
  OAI211_X1 g1075(.A(new_n1275_), .B(new_n954_), .C1(new_n977_), .C2(new_n976_), .ZN(new_n1276_));
  NAND2_X1  g1076(.A1(G390), .A2(new_n978_), .ZN(new_n1277_));
  NAND2_X1  g1077(.A1(new_n1276_), .A2(new_n1277_), .ZN(new_n1278_));
  NAND2_X1  g1078(.A1(G393), .A2(G396), .ZN(new_n1279_));
  NAND2_X1  g1079(.A1(new_n1279_), .A2(new_n1218_), .ZN(new_n1280_));
  XNOR2_X1  g1080(.A(new_n1278_), .B(new_n1280_), .ZN(new_n1281_));
  NAND4_X1  g1081(.A1(new_n1265_), .A2(new_n1267_), .A3(new_n1274_), .A4(new_n1281_), .ZN(new_n1282_));
  INV_X1    g1082(.A(KEYINPUT121), .ZN(new_n1283_));
  NAND2_X1  g1083(.A1(new_n1261_), .A2(new_n1283_), .ZN(new_n1284_));
  NAND4_X1  g1084(.A1(new_n1243_), .A2(new_n1245_), .A3(new_n1253_), .A4(KEYINPUT121), .ZN(new_n1285_));
  NAND2_X1  g1085(.A1(new_n1284_), .A2(new_n1285_), .ZN(new_n1286_));
  INV_X1    g1086(.A(KEYINPUT120), .ZN(new_n1287_));
  NAND4_X1  g1087(.A1(new_n1255_), .A2(new_n1287_), .A3(new_n1258_), .A4(new_n1259_), .ZN(new_n1288_));
  NAND2_X1  g1088(.A1(new_n1258_), .A2(new_n1259_), .ZN(new_n1289_));
  OAI21_X1  g1089(.A(KEYINPUT120), .B1(new_n1246_), .B2(new_n1289_), .ZN(new_n1290_));
  NAND4_X1  g1090(.A1(new_n1274_), .A2(new_n1286_), .A3(new_n1288_), .A4(new_n1290_), .ZN(new_n1291_));
  INV_X1    g1091(.A(KEYINPUT124), .ZN(new_n1292_));
  AND2_X1   g1092(.A1(new_n1276_), .A2(new_n1277_), .ZN(new_n1293_));
  INV_X1    g1093(.A(KEYINPUT123), .ZN(new_n1294_));
  OAI21_X1  g1094(.A(KEYINPUT122), .B1(new_n1280_), .B2(new_n1294_), .ZN(new_n1295_));
  NAND2_X1  g1095(.A1(new_n1293_), .A2(new_n1295_), .ZN(new_n1296_));
  AOI21_X1  g1096(.A(new_n1294_), .B1(new_n1278_), .B2(KEYINPUT122), .ZN(new_n1297_));
  INV_X1    g1097(.A(new_n1280_), .ZN(new_n1298_));
  OAI21_X1  g1098(.A(new_n1296_), .B1(new_n1297_), .B2(new_n1298_), .ZN(new_n1299_));
  INV_X1    g1099(.A(new_n1299_), .ZN(new_n1300_));
  AND3_X1   g1100(.A1(new_n1291_), .A2(new_n1292_), .A3(new_n1300_), .ZN(new_n1301_));
  AOI21_X1  g1101(.A(new_n1292_), .B1(new_n1291_), .B2(new_n1300_), .ZN(new_n1302_));
  OAI21_X1  g1102(.A(new_n1282_), .B1(new_n1301_), .B2(new_n1302_), .ZN(G405));
  XNOR2_X1  g1103(.A(new_n1192_), .B(new_n1222_), .ZN(new_n1304_));
  INV_X1    g1104(.A(new_n1304_), .ZN(new_n1305_));
  OAI21_X1  g1105(.A(KEYINPUT127), .B1(G375), .B2(new_n1222_), .ZN(new_n1306_));
  AND2_X1   g1106(.A1(new_n1306_), .A2(new_n1257_), .ZN(new_n1307_));
  NAND2_X1  g1107(.A1(new_n1299_), .A2(new_n1307_), .ZN(new_n1308_));
  INV_X1    g1108(.A(new_n1308_), .ZN(new_n1309_));
  NOR2_X1   g1109(.A1(new_n1299_), .A2(new_n1307_), .ZN(new_n1310_));
  OAI21_X1  g1110(.A(new_n1305_), .B1(new_n1309_), .B2(new_n1310_), .ZN(new_n1311_));
  OR2_X1    g1111(.A1(new_n1299_), .A2(new_n1307_), .ZN(new_n1312_));
  NAND3_X1  g1112(.A1(new_n1312_), .A2(new_n1304_), .A3(new_n1308_), .ZN(new_n1313_));
  NAND2_X1  g1113(.A1(new_n1311_), .A2(new_n1313_), .ZN(G402));
endmodule


