//Secret key is'1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_c7552" written by ABC on Wed Oct 26 14:18:04 2022

module locked_c7552 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G5, G9, G12, G15,
    G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55,
    G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87,
    G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113,
    G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141,
    G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159,
    G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171,
    G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183,
    G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195,
    G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207,
    G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219,
    G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231,
    G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197,
    G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208,
    G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698,
    G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393,
    G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526,
    G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G5, G9,
    G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53,
    G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69,
    G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85,
    G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112,
    G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138,
    G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218,
    G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230,
    G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339,
    G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204,
    G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256,
    G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749,
    G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437,
    G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_n426_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1114_, new_n1115_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1128_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1305_, new_n1307_, new_n1308_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1339_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1354_,
    new_n1355_, new_n1358_, new_n1359_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1382_, new_n1383_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1414_, new_n1415_, new_n1416_,
    new_n1419_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1433_, new_n1434_, new_n1435_, new_n1438_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_;
  BUF_X1    g0000(.A(G1), .Z(G2));
  BUF_X1    g0001(.A(G1), .Z(G3));
  BUF_X1    g0002(.A(G1459), .Z(G450));
  BUF_X1    g0003(.A(G1469), .Z(G448));
  BUF_X1    g0004(.A(G1480), .Z(G444));
  BUF_X1    g0005(.A(G1486), .Z(G442));
  BUF_X1    g0006(.A(G1492), .Z(G440));
  BUF_X1    g0007(.A(G1496), .Z(G438));
  BUF_X1    g0008(.A(G2208), .Z(G496));
  BUF_X1    g0009(.A(G2218), .Z(G494));
  BUF_X1    g0010(.A(G2224), .Z(G492));
  XNOR2_X1  g0011(.A(KEYINPUT0), .B(G2230), .ZN(G490));
  BUF_X1    g0012(.A(G2236), .Z(G488));
  BUF_X1    g0013(.A(G2239), .Z(G486));
  BUF_X1    g0014(.A(G2247), .Z(G484));
  BUF_X1    g0015(.A(G2253), .Z(G482));
  BUF_X1    g0016(.A(G2256), .Z(G480));
  BUF_X1    g0017(.A(G3698), .Z(G560));
  BUF_X1    g0018(.A(G3701), .Z(G542));
  BUF_X1    g0019(.A(G3705), .Z(G558));
  BUF_X1    g0020(.A(G3711), .Z(G556));
  BUF_X1    g0021(.A(G3717), .Z(G554));
  BUF_X1    g0022(.A(G3723), .Z(G552));
  BUF_X1    g0023(.A(G3729), .Z(G550));
  BUF_X1    g0024(.A(G3737), .Z(G548));
  BUF_X1    g0025(.A(G3743), .Z(G546));
  BUF_X1    g0026(.A(G3749), .Z(G544));
  BUF_X1    g0027(.A(G4393), .Z(G540));
  XNOR2_X1  g0028(.A(KEYINPUT1), .B(G4400), .ZN(G538));
  BUF_X1    g0029(.A(G4405), .Z(G536));
  BUF_X1    g0030(.A(G4410), .Z(G534));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G4415), .Z(G532));
  BUF_X1    g0032(.A(G4420), .Z(G530));
  BUF_X1    g0033(.A(G4427), .Z(G528));
  BUF_X1    g0034(.A(G4432), .Z(G526));
  BUF_X1    g0035(.A(G4437), .Z(G524));
  INV_X1    g0036(.A(G15), .ZN(G279));
  BUF_X1    g0037(.A(G1462), .Z(G436));
  BUF_X1    g0038(.A(G2211), .Z(G478));
  BUF_X1    g0039(.A(G4394), .Z(G522));
  OR2_X1    g0040(.A1(G5), .A2(G57), .ZN(G402));
  NAND4_X1  g0041(.A1(G150), .A2(G184), .A3(G228), .A4(G240), .ZN(G404));
  NAND4_X1  g0042(.A1(G152), .A2(G210), .A3(G218), .A4(G230), .ZN(G406));
  NAND4_X1  g0043(.A1(G182), .A2(G183), .A3(G185), .A4(G186), .ZN(G408));
  NAND4_X1  g0044(.A1(G162), .A2(G172), .A3(G188), .A4(G199), .ZN(G410));
  BUF_X1    g0045(.A(G1), .Z(G432));
  BUF_X1    g0046(.A(G106), .Z(G446));
  INV_X1    g0047(.A(G5), .ZN(new_n426_));
  NAND2_X1  g0048(.A1(new_n426_), .A2(G1197), .ZN(G284));
  INV_X1    g0049(.A(G15), .ZN(G286));
  NAND2_X1  g0050(.A1(new_n426_), .A2(G1197), .ZN(G289));
  NAND3_X1  g0051(.A1(new_n426_), .A2(G133), .A3(G134), .ZN(G292));
  INV_X1    g0052(.A(G15), .ZN(G341));
  NAND3_X1  g0053(.A1(new_n426_), .A2(G133), .A3(G134), .ZN(G281));
  BUF_X1    g0054(.A(G1), .Z(G453));
  AND2_X1   g0055(.A1(G1), .A2(G163), .ZN(G278));
  INV_X1    g0056(.A(G41), .ZN(new_n435_));
  OR3_X1    g0057(.A1(new_n435_), .A2(G18), .A3(G3701), .ZN(new_n436_));
  INV_X1    g0058(.A(G18), .ZN(new_n437_));
  NAND3_X1  g0059(.A1(new_n437_), .A2(new_n435_), .A3(G3701), .ZN(new_n438_));
  NAND2_X1  g0060(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g0061(.A(new_n439_), .B(G4526), .ZN(new_n440_));
  XNOR2_X1  g0062(.A(new_n440_), .B(KEYINPUT3), .ZN(G373));
  NAND2_X1  g0063(.A1(G1496), .A2(G4528), .ZN(new_n442_));
  INV_X1    g0064(.A(G1492), .ZN(new_n443_));
  NOR2_X1   g0065(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g0066(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g0067(.A1(new_n445_), .A2(G38), .ZN(new_n446_));
  NAND2_X1  g0068(.A1(G9), .A2(G12), .ZN(new_n447_));
  OAI21_X1  g0069(.A(new_n447_), .B1(new_n437_), .B2(G215), .ZN(new_n448_));
  NAND2_X1  g0070(.A1(new_n448_), .A2(G106), .ZN(new_n449_));
  INV_X1    g0071(.A(G106), .ZN(new_n450_));
  OAI211_X1 g0072(.A(new_n447_), .B(new_n450_), .C1(new_n437_), .C2(G215), .ZN(new_n451_));
  AND2_X1   g0073(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g0074(.A(G216), .ZN(new_n453_));
  NAND2_X1  g0075(.A1(new_n453_), .A2(G18), .ZN(new_n454_));
  INV_X1    g0076(.A(G1469), .ZN(new_n455_));
  NAND3_X1  g0077(.A1(new_n454_), .A2(new_n455_), .A3(new_n447_), .ZN(new_n456_));
  INV_X1    g0078(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g0079(.A(new_n455_), .B1(new_n454_), .B2(new_n447_), .ZN(new_n458_));
  NOR2_X1   g0080(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g0081(.A1(new_n452_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g0082(.A(G1486), .ZN(new_n461_));
  OR2_X1    g0083(.A1(new_n437_), .A2(G213), .ZN(new_n462_));
  AOI21_X1  g0084(.A(new_n461_), .B1(new_n462_), .B2(new_n447_), .ZN(new_n463_));
  INV_X1    g0085(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g0086(.A1(new_n462_), .A2(new_n461_), .A3(new_n447_), .ZN(new_n465_));
  NAND2_X1  g0087(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g0088(.A(G1480), .ZN(new_n467_));
  INV_X1    g0089(.A(G214), .ZN(new_n468_));
  NAND2_X1  g0090(.A1(new_n468_), .A2(G18), .ZN(new_n469_));
  AOI21_X1  g0091(.A(new_n467_), .B1(new_n469_), .B2(new_n447_), .ZN(new_n470_));
  INV_X1    g0092(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g0093(.A1(new_n469_), .A2(new_n467_), .A3(new_n447_), .ZN(new_n472_));
  NAND2_X1  g0094(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g0095(.A(G209), .ZN(new_n474_));
  NAND2_X1  g0096(.A1(new_n474_), .A2(G18), .ZN(new_n475_));
  INV_X1    g0097(.A(G1462), .ZN(new_n476_));
  NAND3_X1  g0098(.A1(new_n475_), .A2(new_n476_), .A3(new_n447_), .ZN(new_n477_));
  NOR3_X1   g0099(.A1(new_n466_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g0100(.A(KEYINPUT18), .ZN(new_n479_));
  AOI21_X1  g0101(.A(new_n460_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g0102(.A(new_n480_), .B1(new_n479_), .B2(new_n478_), .ZN(new_n481_));
  AND2_X1   g0103(.A1(new_n472_), .A2(new_n451_), .ZN(new_n482_));
  NAND2_X1  g0104(.A1(new_n449_), .A2(new_n451_), .ZN(new_n483_));
  OAI21_X1  g0105(.A(new_n482_), .B1(new_n483_), .B2(new_n456_), .ZN(new_n484_));
  NAND3_X1  g0106(.A1(new_n484_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n485_));
  NAND3_X1  g0107(.A1(new_n481_), .A2(new_n465_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g0108(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g0109(.A(G4528), .ZN(new_n488_));
  NOR3_X1   g0110(.A1(new_n443_), .A2(new_n488_), .A3(G38), .ZN(new_n489_));
  INV_X1    g0111(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g0112(.A(G38), .B1(new_n443_), .B2(new_n488_), .ZN(new_n491_));
  NAND2_X1  g0113(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g0114(.A(new_n442_), .B(G38), .ZN(new_n493_));
  OR2_X1    g0115(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g0116(.A(new_n446_), .B1(new_n487_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g0117(.A(new_n447_), .B1(new_n437_), .B2(G153), .ZN(new_n496_));
  XNOR2_X1  g0118(.A(new_n496_), .B(KEYINPUT6), .ZN(new_n497_));
  OR2_X1    g0119(.A1(new_n497_), .A2(G2256), .ZN(new_n498_));
  INV_X1    g0120(.A(G154), .ZN(new_n499_));
  AOI21_X1  g0121(.A(new_n437_), .B1(KEYINPUT5), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g0122(.A(new_n500_), .B1(KEYINPUT5), .B2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g0123(.A1(new_n501_), .A2(new_n447_), .ZN(new_n502_));
  NAND2_X1  g0124(.A1(new_n502_), .A2(G2253), .ZN(new_n503_));
  INV_X1    g0125(.A(new_n503_), .ZN(new_n504_));
  OR2_X1    g0126(.A1(new_n437_), .A2(G155), .ZN(new_n505_));
  AND2_X1   g0127(.A1(new_n505_), .A2(new_n447_), .ZN(new_n506_));
  INV_X1    g0128(.A(G2247), .ZN(new_n507_));
  OR2_X1    g0129(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g0130(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  INV_X1    g0131(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g0132(.A(new_n447_), .ZN(new_n511_));
  INV_X1    g0133(.A(G156), .ZN(new_n512_));
  AOI21_X1  g0134(.A(new_n511_), .B1(G18), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g0135(.A(G2239), .ZN(new_n514_));
  NAND2_X1  g0136(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g0137(.A(new_n515_), .ZN(new_n516_));
  OAI21_X1  g0138(.A(new_n508_), .B1(new_n510_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g0139(.A(new_n502_), .ZN(new_n518_));
  INV_X1    g0140(.A(G2253), .ZN(new_n519_));
  NAND2_X1  g0141(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g0142(.A(new_n504_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g0143(.A1(new_n497_), .A2(G2256), .ZN(new_n522_));
  NAND2_X1  g0144(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g0145(.A(G135), .ZN(new_n524_));
  NOR2_X1   g0146(.A1(new_n524_), .A2(G18), .ZN(new_n525_));
  AOI21_X1  g0147(.A(new_n525_), .B1(G18), .B2(G158), .ZN(new_n526_));
  OR2_X1    g0148(.A1(new_n526_), .A2(G2230), .ZN(new_n527_));
  INV_X1    g0149(.A(KEYINPUT8), .ZN(new_n528_));
  INV_X1    g0150(.A(G144), .ZN(new_n529_));
  AOI21_X1  g0151(.A(G18), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g0152(.A(new_n530_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n531_));
  NAND2_X1  g0153(.A1(G18), .A2(G159), .ZN(new_n532_));
  NAND2_X1  g0154(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g0155(.A(G2224), .ZN(new_n534_));
  NAND2_X1  g0156(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g0157(.A1(new_n526_), .A2(G2230), .ZN(new_n536_));
  INV_X1    g0158(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g0159(.A(new_n527_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g0160(.A1(new_n531_), .A2(G2224), .A3(new_n532_), .ZN(new_n539_));
  NAND2_X1  g0161(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g0162(.A1(new_n527_), .A2(new_n536_), .ZN(new_n541_));
  NOR2_X1   g0163(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g0164(.A1(G18), .A2(G160), .ZN(new_n543_));
  INV_X1    g0165(.A(G138), .ZN(new_n544_));
  OAI21_X1  g0166(.A(new_n543_), .B1(new_n544_), .B2(G18), .ZN(new_n545_));
  INV_X1    g0167(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g0168(.A(G2218), .ZN(new_n547_));
  NAND2_X1  g0169(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g0170(.A(KEYINPUT9), .ZN(new_n549_));
  NAND2_X1  g0171(.A1(new_n545_), .A2(G2218), .ZN(new_n550_));
  NAND3_X1  g0172(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g0173(.A(new_n550_), .ZN(new_n552_));
  NAND2_X1  g0174(.A1(new_n552_), .A2(KEYINPUT9), .ZN(new_n553_));
  NAND2_X1  g0175(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g0176(.A1(new_n437_), .A2(G147), .ZN(new_n555_));
  INV_X1    g0177(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g0178(.A(new_n556_), .B1(G18), .B2(G151), .ZN(new_n557_));
  NOR2_X1   g0179(.A1(new_n557_), .A2(G2211), .ZN(new_n558_));
  INV_X1    g0180(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g0181(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g0182(.A(new_n538_), .B1(new_n542_), .B2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g0183(.A1(new_n546_), .A2(G2218), .ZN(new_n562_));
  NAND2_X1  g0184(.A1(new_n542_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g0185(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g0186(.A(new_n447_), .B1(new_n437_), .B2(G157), .ZN(new_n565_));
  XNOR2_X1  g0187(.A(new_n565_), .B(KEYINPUT7), .ZN(new_n566_));
  INV_X1    g0188(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g0189(.A1(new_n567_), .A2(G2236), .ZN(new_n568_));
  NAND2_X1  g0190(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  OR2_X1    g0191(.A1(new_n567_), .A2(G2236), .ZN(new_n570_));
  NAND2_X1  g0192(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g0193(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g0194(.A(new_n508_), .ZN(new_n573_));
  NOR2_X1   g0195(.A1(new_n573_), .A2(new_n510_), .ZN(new_n574_));
  NAND3_X1  g0196(.A1(new_n574_), .A2(new_n520_), .A3(new_n503_), .ZN(new_n575_));
  NOR2_X1   g0197(.A1(new_n513_), .A2(new_n514_), .ZN(new_n576_));
  NOR2_X1   g0198(.A1(new_n516_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g0199(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g0200(.A1(new_n498_), .A2(new_n522_), .ZN(new_n579_));
  NOR3_X1   g0201(.A1(new_n575_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g0202(.A(new_n580_), .ZN(new_n581_));
  OAI211_X1 g0203(.A(new_n498_), .B(new_n523_), .C1(new_n572_), .C2(new_n581_), .ZN(new_n582_));
  INV_X1    g0204(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g0205(.A1(new_n557_), .A2(G2211), .ZN(new_n584_));
  INV_X1    g0206(.A(new_n584_), .ZN(new_n585_));
  NOR3_X1   g0207(.A1(new_n554_), .A2(new_n585_), .A3(new_n558_), .ZN(new_n586_));
  NAND2_X1  g0208(.A1(new_n586_), .A2(new_n542_), .ZN(new_n587_));
  NAND2_X1  g0209(.A1(new_n570_), .A2(new_n568_), .ZN(new_n588_));
  OR2_X1    g0210(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g0211(.A(new_n589_), .B(KEYINPUT10), .Z(new_n590_));
  NAND2_X1  g0212(.A1(new_n590_), .A2(new_n580_), .ZN(new_n591_));
  NAND2_X1  g0213(.A1(new_n437_), .A2(G130), .ZN(new_n592_));
  INV_X1    g0214(.A(G234), .ZN(new_n593_));
  OAI21_X1  g0215(.A(new_n592_), .B1(new_n437_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g0216(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g0217(.A1(new_n595_), .A2(G3729), .ZN(new_n596_));
  INV_X1    g0218(.A(G3729), .ZN(new_n597_));
  NAND2_X1  g0219(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g0220(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g0221(.A(new_n599_), .B(KEYINPUT13), .ZN(new_n600_));
  NAND2_X1  g0222(.A1(new_n437_), .A2(G127), .ZN(new_n601_));
  NAND2_X1  g0223(.A1(G18), .A2(G233), .ZN(new_n602_));
  AND2_X1   g0224(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g0225(.A1(new_n603_), .A2(G3737), .ZN(new_n604_));
  NAND2_X1  g0226(.A1(new_n603_), .A2(G3737), .ZN(new_n605_));
  INV_X1    g0227(.A(new_n605_), .ZN(new_n606_));
  NOR3_X1   g0228(.A1(new_n600_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g0229(.A1(new_n437_), .A2(G124), .ZN(new_n608_));
  INV_X1    g0230(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g0231(.A(new_n609_), .B1(G18), .B2(G232), .ZN(new_n610_));
  OR2_X1    g0232(.A1(new_n610_), .A2(G3743), .ZN(new_n611_));
  NAND2_X1  g0233(.A1(new_n610_), .A2(G3743), .ZN(new_n612_));
  NAND2_X1  g0234(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g0235(.A1(new_n437_), .A2(G100), .ZN(new_n614_));
  AOI21_X1  g0236(.A(new_n614_), .B1(G18), .B2(G231), .ZN(new_n615_));
  OR2_X1    g0237(.A1(new_n615_), .A2(G3749), .ZN(new_n616_));
  NAND2_X1  g0238(.A1(new_n615_), .A2(G3749), .ZN(new_n617_));
  NAND2_X1  g0239(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g0240(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g0241(.A1(new_n607_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g0242(.A(G235), .ZN(new_n621_));
  NOR2_X1   g0243(.A1(new_n621_), .A2(KEYINPUT12), .ZN(new_n622_));
  INV_X1    g0244(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g0245(.A(new_n437_), .B1(KEYINPUT12), .B2(new_n621_), .ZN(new_n624_));
  AOI22_X1  g0246(.A1(new_n623_), .A2(new_n624_), .B1(new_n437_), .B2(G103), .ZN(new_n625_));
  OR2_X1    g0247(.A1(new_n625_), .A2(G3723), .ZN(new_n626_));
  NAND2_X1  g0248(.A1(new_n625_), .A2(G3723), .ZN(new_n627_));
  NAND2_X1  g0249(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g0250(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g0251(.A1(G18), .A2(G237), .ZN(new_n630_));
  INV_X1    g0252(.A(G26), .ZN(new_n631_));
  OAI21_X1  g0253(.A(new_n630_), .B1(new_n631_), .B2(G18), .ZN(new_n632_));
  INV_X1    g0254(.A(G3711), .ZN(new_n633_));
  NAND2_X1  g0255(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g0256(.A(KEYINPUT11), .B(G3711), .ZN(new_n635_));
  OAI21_X1  g0257(.A(new_n634_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g0258(.A1(G18), .A2(G236), .ZN(new_n637_));
  INV_X1    g0259(.A(G23), .ZN(new_n638_));
  OAI21_X1  g0260(.A(new_n637_), .B1(new_n638_), .B2(G18), .ZN(new_n639_));
  INV_X1    g0261(.A(G3717), .ZN(new_n640_));
  NAND2_X1  g0262(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g0263(.A(new_n637_), .B(G3717), .C1(G18), .C2(new_n638_), .ZN(new_n642_));
  NAND2_X1  g0264(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g0265(.A1(new_n636_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g0266(.A1(G18), .A2(G238), .ZN(new_n645_));
  INV_X1    g0267(.A(G29), .ZN(new_n646_));
  OAI21_X1  g0268(.A(new_n645_), .B1(new_n646_), .B2(G18), .ZN(new_n647_));
  INV_X1    g0269(.A(G3705), .ZN(new_n648_));
  NAND2_X1  g0270(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g0271(.A(new_n645_), .B(G3705), .C1(G18), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g0272(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g0273(.A1(new_n651_), .A2(new_n439_), .ZN(new_n652_));
  NAND4_X1  g0274(.A1(new_n629_), .A2(G4526), .A3(new_n644_), .A4(new_n652_), .ZN(new_n653_));
  NOR2_X1   g0275(.A1(new_n620_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g0276(.A(KEYINPUT17), .ZN(new_n655_));
  NAND2_X1  g0277(.A1(new_n437_), .A2(G32), .ZN(new_n656_));
  NAND2_X1  g0278(.A1(G18), .A2(G221), .ZN(new_n657_));
  NAND2_X1  g0279(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g0280(.A(KEYINPUT15), .ZN(new_n659_));
  NAND2_X1  g0281(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g0282(.A1(new_n656_), .A2(KEYINPUT15), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g0283(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g0284(.A(G4427), .ZN(new_n663_));
  NAND2_X1  g0285(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g0286(.A1(new_n660_), .A2(G4427), .A3(new_n661_), .ZN(new_n665_));
  AOI21_X1  g0287(.A(KEYINPUT16), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g0288(.A1(new_n662_), .A2(KEYINPUT16), .A3(G4427), .ZN(new_n667_));
  INV_X1    g0289(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g0290(.A(new_n655_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g0291(.A(KEYINPUT16), .ZN(new_n670_));
  INV_X1    g0292(.A(new_n665_), .ZN(new_n671_));
  AOI21_X1  g0293(.A(G4427), .B1(new_n660_), .B2(new_n661_), .ZN(new_n672_));
  OAI21_X1  g0294(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g0295(.A1(new_n673_), .A2(KEYINPUT17), .A3(new_n667_), .ZN(new_n674_));
  NAND2_X1  g0296(.A1(new_n669_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g0297(.A1(new_n437_), .A2(G35), .ZN(new_n676_));
  INV_X1    g0298(.A(G222), .ZN(new_n677_));
  OAI21_X1  g0299(.A(new_n676_), .B1(new_n437_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g0300(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g0301(.A1(new_n679_), .A2(G4420), .ZN(new_n680_));
  INV_X1    g0302(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g0303(.A1(new_n679_), .A2(G4420), .ZN(new_n682_));
  NOR2_X1   g0304(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g0305(.A1(new_n437_), .A2(G50), .ZN(new_n684_));
  INV_X1    g0306(.A(G220), .ZN(new_n685_));
  OAI21_X1  g0307(.A(new_n684_), .B1(new_n437_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g0308(.A(new_n686_), .ZN(new_n687_));
  OR2_X1    g0309(.A1(new_n687_), .A2(G4432), .ZN(new_n688_));
  NAND2_X1  g0310(.A1(new_n687_), .A2(G4432), .ZN(new_n689_));
  NAND2_X1  g0311(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g0312(.A1(new_n437_), .A2(G66), .ZN(new_n691_));
  INV_X1    g0313(.A(G219), .ZN(new_n692_));
  OAI21_X1  g0314(.A(new_n691_), .B1(new_n437_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g0315(.A(G4437), .ZN(new_n694_));
  XNOR2_X1  g0316(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NOR2_X1   g0317(.A1(new_n690_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g0318(.A1(G18), .A2(G226), .ZN(new_n697_));
  INV_X1    g0319(.A(G97), .ZN(new_n698_));
  OAI21_X1  g0320(.A(new_n697_), .B1(new_n698_), .B2(G18), .ZN(new_n699_));
  INV_X1    g0321(.A(G4400), .ZN(new_n700_));
  NAND2_X1  g0322(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g0323(.A1(new_n437_), .A2(G97), .ZN(new_n702_));
  NAND3_X1  g0324(.A1(new_n702_), .A2(G4400), .A3(new_n697_), .ZN(new_n703_));
  AND2_X1   g0325(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g0326(.A1(new_n437_), .A2(G118), .ZN(new_n705_));
  NAND2_X1  g0327(.A1(G18), .A2(G217), .ZN(new_n706_));
  NAND3_X1  g0328(.A1(new_n705_), .A2(G4394), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g0329(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g0330(.A(G4394), .B1(new_n705_), .B2(new_n706_), .ZN(new_n709_));
  NOR2_X1   g0331(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g0332(.A1(new_n437_), .A2(G121), .ZN(new_n711_));
  NAND2_X1  g0333(.A1(G18), .A2(G224), .ZN(new_n712_));
  NAND3_X1  g0334(.A1(new_n711_), .A2(G4410), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g0335(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g0336(.A(G4410), .B1(new_n711_), .B2(new_n712_), .ZN(new_n715_));
  NOR2_X1   g0337(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g0338(.A1(G18), .A2(G225), .ZN(new_n717_));
  INV_X1    g0339(.A(G94), .ZN(new_n718_));
  OAI211_X1 g0340(.A(new_n717_), .B(G4405), .C1(G18), .C2(new_n718_), .ZN(new_n719_));
  INV_X1    g0341(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g0342(.A1(new_n437_), .A2(G94), .ZN(new_n721_));
  AOI21_X1  g0343(.A(G4405), .B1(new_n721_), .B2(new_n717_), .ZN(new_n722_));
  NOR2_X1   g0344(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND4_X1  g0345(.A1(new_n704_), .A2(new_n710_), .A3(new_n716_), .A4(new_n723_), .ZN(new_n724_));
  MUX2_X1   g0346(.A(G47), .B(G223), .S(G18), .Z(new_n725_));
  INV_X1    g0347(.A(G4415), .ZN(new_n726_));
  OR2_X1    g0348(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g0349(.A1(new_n725_), .A2(new_n726_), .ZN(new_n728_));
  NAND2_X1  g0350(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g0351(.A1(new_n724_), .A2(new_n729_), .ZN(new_n730_));
  AND4_X1   g0352(.A1(new_n675_), .A2(new_n683_), .A3(new_n696_), .A4(new_n730_), .ZN(new_n731_));
  NAND2_X1  g0353(.A1(new_n654_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g0354(.A(new_n583_), .B1(new_n591_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g0355(.A(KEYINPUT4), .B1(new_n475_), .B2(new_n447_), .ZN(new_n734_));
  INV_X1    g0356(.A(new_n734_), .ZN(new_n735_));
  OAI211_X1 g0357(.A(new_n447_), .B(KEYINPUT4), .C1(new_n437_), .C2(G209), .ZN(new_n736_));
  NAND3_X1  g0358(.A1(new_n735_), .A2(G1462), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g0359(.A(new_n736_), .ZN(new_n738_));
  OAI21_X1  g0360(.A(new_n476_), .B1(new_n738_), .B2(new_n734_), .ZN(new_n739_));
  NAND3_X1  g0361(.A1(new_n737_), .A2(new_n739_), .A3(new_n459_), .ZN(new_n740_));
  NOR2_X1   g0362(.A1(new_n473_), .A2(new_n483_), .ZN(new_n741_));
  INV_X1    g0363(.A(new_n741_), .ZN(new_n742_));
  NOR4_X1   g0364(.A1(new_n740_), .A2(new_n494_), .A3(new_n742_), .A4(new_n466_), .ZN(new_n743_));
  AOI21_X1  g0365(.A(new_n495_), .B1(new_n733_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g0366(.A1(new_n611_), .A2(new_n616_), .ZN(new_n745_));
  AND2_X1   g0367(.A1(new_n745_), .A2(new_n617_), .ZN(new_n746_));
  XNOR2_X1  g0368(.A(new_n598_), .B(KEYINPUT14), .ZN(new_n747_));
  INV_X1    g0369(.A(new_n604_), .ZN(new_n748_));
  AOI21_X1  g0370(.A(new_n606_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g0371(.A(new_n746_), .B1(new_n749_), .B2(new_n619_), .ZN(new_n750_));
  INV_X1    g0372(.A(new_n626_), .ZN(new_n751_));
  INV_X1    g0373(.A(new_n643_), .ZN(new_n752_));
  NAND2_X1  g0374(.A1(new_n437_), .A2(G26), .ZN(new_n753_));
  AOI21_X1  g0375(.A(G3711), .B1(new_n753_), .B2(new_n630_), .ZN(new_n754_));
  INV_X1    g0376(.A(new_n632_), .ZN(new_n755_));
  XOR2_X1   g0377(.A(KEYINPUT11), .B(G3711), .Z(new_n756_));
  AOI21_X1  g0378(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g0379(.A1(new_n437_), .A2(G29), .ZN(new_n758_));
  AOI21_X1  g0380(.A(G3705), .B1(new_n758_), .B2(new_n645_), .ZN(new_n759_));
  NAND3_X1  g0381(.A1(new_n752_), .A2(new_n757_), .A3(new_n759_), .ZN(new_n760_));
  AND2_X1   g0382(.A1(new_n635_), .A2(new_n632_), .ZN(new_n761_));
  NOR3_X1   g0383(.A1(new_n435_), .A2(G18), .A3(G3701), .ZN(new_n762_));
  AND3_X1   g0384(.A1(new_n649_), .A2(new_n762_), .A3(new_n650_), .ZN(new_n763_));
  AOI21_X1  g0385(.A(new_n761_), .B1(new_n763_), .B2(new_n757_), .ZN(new_n764_));
  INV_X1    g0386(.A(new_n642_), .ZN(new_n765_));
  OAI211_X1 g0387(.A(new_n641_), .B(new_n760_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g0388(.A(new_n751_), .B1(new_n766_), .B2(new_n627_), .ZN(new_n767_));
  OAI21_X1  g0389(.A(new_n750_), .B1(new_n620_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g0390(.A1(new_n768_), .A2(new_n731_), .ZN(new_n769_));
  INV_X1    g0391(.A(new_n682_), .ZN(new_n770_));
  NAND2_X1  g0392(.A1(new_n770_), .A2(new_n664_), .ZN(new_n771_));
  OAI211_X1 g0393(.A(new_n771_), .B(new_n689_), .C1(new_n675_), .C2(new_n672_), .ZN(new_n772_));
  NAND2_X1  g0394(.A1(new_n772_), .A2(new_n688_), .ZN(new_n773_));
  INV_X1    g0395(.A(new_n695_), .ZN(new_n774_));
  NAND2_X1  g0396(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AND3_X1   g0397(.A1(new_n675_), .A2(new_n683_), .A3(new_n696_), .ZN(new_n776_));
  INV_X1    g0398(.A(G121), .ZN(new_n777_));
  OAI21_X1  g0399(.A(new_n712_), .B1(new_n777_), .B2(G18), .ZN(new_n778_));
  INV_X1    g0400(.A(G4410), .ZN(new_n779_));
  NAND2_X1  g0401(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OR3_X1    g0402(.A1(new_n729_), .A2(KEYINPUT19), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g0403(.A(KEYINPUT19), .B1(new_n729_), .B2(new_n780_), .ZN(new_n782_));
  NAND3_X1  g0404(.A1(new_n716_), .A2(new_n727_), .A3(new_n722_), .ZN(new_n783_));
  NAND4_X1  g0405(.A1(new_n781_), .A2(new_n728_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n784_));
  INV_X1    g0406(.A(new_n729_), .ZN(new_n785_));
  OAI21_X1  g0407(.A(new_n717_), .B1(new_n718_), .B2(G18), .ZN(new_n786_));
  INV_X1    g0408(.A(G4405), .ZN(new_n787_));
  NAND2_X1  g0409(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g0410(.A1(new_n780_), .A2(new_n788_), .A3(new_n713_), .A4(new_n719_), .ZN(new_n789_));
  INV_X1    g0411(.A(new_n789_), .ZN(new_n790_));
  NAND3_X1  g0412(.A1(new_n701_), .A2(new_n703_), .A3(new_n709_), .ZN(new_n791_));
  NAND2_X1  g0413(.A1(new_n791_), .A2(new_n701_), .ZN(new_n792_));
  AND3_X1   g0414(.A1(new_n785_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  OR2_X1    g0415(.A1(new_n784_), .A2(new_n793_), .ZN(new_n794_));
  AOI22_X1  g0416(.A1(new_n776_), .A2(new_n794_), .B1(new_n694_), .B2(new_n693_), .ZN(new_n795_));
  NAND3_X1  g0417(.A1(new_n769_), .A2(new_n775_), .A3(new_n795_), .ZN(new_n796_));
  AND3_X1   g0418(.A1(new_n796_), .A2(new_n590_), .A3(new_n580_), .ZN(new_n797_));
  NAND2_X1  g0419(.A1(new_n797_), .A2(new_n743_), .ZN(new_n798_));
  NAND2_X1  g0420(.A1(new_n744_), .A2(new_n798_), .ZN(G246));
  NOR2_X1   g0421(.A1(new_n488_), .A2(G2204), .ZN(new_n800_));
  XNOR2_X1  g0422(.A(new_n800_), .B(KEYINPUT24), .ZN(new_n801_));
  OR2_X1    g0423(.A1(new_n488_), .A2(G1455), .ZN(new_n802_));
  OAI21_X1  g0424(.A(G38), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g0425(.A(new_n447_), .B1(new_n437_), .B2(G166), .ZN(new_n804_));
  NAND2_X1  g0426(.A1(G18), .A2(G1486), .ZN(new_n805_));
  OAI21_X1  g0427(.A(new_n805_), .B1(G18), .B2(G88), .ZN(new_n806_));
  XNOR2_X1  g0428(.A(new_n804_), .B(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g0429(.A(new_n807_), .B(KEYINPUT22), .ZN(new_n808_));
  NOR2_X1   g0430(.A1(G18), .A2(G112), .ZN(new_n809_));
  AOI21_X1  g0431(.A(new_n809_), .B1(G18), .B2(G1480), .ZN(new_n810_));
  INV_X1    g0432(.A(new_n810_), .ZN(new_n811_));
  OAI21_X1  g0433(.A(new_n447_), .B1(new_n437_), .B2(G167), .ZN(new_n812_));
  AND2_X1   g0434(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OR2_X1    g0435(.A1(new_n808_), .A2(new_n813_), .ZN(new_n814_));
  OR2_X1    g0436(.A1(new_n437_), .A2(G168), .ZN(new_n815_));
  NAND2_X1  g0437(.A1(new_n815_), .A2(new_n447_), .ZN(new_n816_));
  NAND2_X1  g0438(.A1(G18), .A2(G106), .ZN(new_n817_));
  OAI21_X1  g0439(.A(new_n817_), .B1(G18), .B2(G87), .ZN(new_n818_));
  NOR2_X1   g0440(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g0441(.A1(new_n811_), .A2(new_n812_), .ZN(new_n820_));
  NAND2_X1  g0442(.A1(G18), .A2(G1462), .ZN(new_n821_));
  OAI21_X1  g0443(.A(new_n821_), .B1(G18), .B2(G113), .ZN(new_n822_));
  NAND2_X1  g0444(.A1(G18), .A2(G1469), .ZN(new_n823_));
  OAI21_X1  g0445(.A(new_n823_), .B1(G18), .B2(G111), .ZN(new_n824_));
  NOR2_X1   g0446(.A1(new_n437_), .A2(G169), .ZN(new_n825_));
  OAI21_X1  g0447(.A(new_n822_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g0448(.A1(new_n826_), .A2(new_n447_), .ZN(new_n827_));
  INV_X1    g0449(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g0450(.A(new_n447_), .B1(new_n437_), .B2(G169), .ZN(new_n829_));
  AOI22_X1  g0451(.A1(new_n816_), .A2(new_n818_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n830_));
  AOI211_X1 g0452(.A(new_n819_), .B(new_n820_), .C1(new_n828_), .C2(new_n830_), .ZN(new_n831_));
  OAI22_X1  g0453(.A1(new_n814_), .A2(new_n831_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n832_));
  OAI21_X1  g0454(.A(new_n447_), .B1(new_n437_), .B2(G174), .ZN(new_n833_));
  INV_X1    g0455(.A(new_n833_), .ZN(new_n834_));
  NOR2_X1   g0456(.A1(G18), .A2(G109), .ZN(new_n835_));
  AOI21_X1  g0457(.A(new_n835_), .B1(G18), .B2(G2253), .ZN(new_n836_));
  NOR2_X1   g0458(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g0459(.A(new_n837_), .ZN(new_n838_));
  NOR2_X1   g0460(.A1(G18), .A2(G86), .ZN(new_n839_));
  AOI21_X1  g0461(.A(new_n839_), .B1(G18), .B2(G2247), .ZN(new_n840_));
  OR2_X1    g0462(.A1(new_n437_), .A2(G175), .ZN(new_n841_));
  NAND3_X1  g0463(.A1(new_n840_), .A2(new_n447_), .A3(new_n841_), .ZN(new_n842_));
  NOR2_X1   g0464(.A1(new_n437_), .A2(G173), .ZN(new_n843_));
  NOR2_X1   g0465(.A1(new_n843_), .A2(new_n511_), .ZN(new_n844_));
  INV_X1    g0466(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g0467(.A1(G18), .A2(G2256), .ZN(new_n846_));
  OAI21_X1  g0468(.A(new_n846_), .B1(G18), .B2(G110), .ZN(new_n847_));
  NAND2_X1  g0469(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g0470(.A(new_n840_), .ZN(new_n849_));
  NAND2_X1  g0471(.A1(new_n841_), .A2(new_n447_), .ZN(new_n850_));
  NAND2_X1  g0472(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g0473(.A1(new_n838_), .A2(new_n842_), .A3(new_n848_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g0474(.A(new_n836_), .ZN(new_n853_));
  OAI22_X1  g0475(.A1(new_n845_), .A2(new_n847_), .B1(new_n853_), .B2(new_n833_), .ZN(new_n854_));
  NOR2_X1   g0476(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g0477(.A(new_n447_), .B1(new_n437_), .B2(G176), .ZN(new_n856_));
  NAND2_X1  g0478(.A1(G18), .A2(G2239), .ZN(new_n857_));
  OAI21_X1  g0479(.A(new_n857_), .B1(G18), .B2(G63), .ZN(new_n858_));
  NOR2_X1   g0480(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g0481(.A1(new_n855_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g0482(.A1(new_n837_), .A2(new_n842_), .ZN(new_n861_));
  OAI21_X1  g0483(.A(new_n848_), .B1(new_n861_), .B2(new_n854_), .ZN(new_n862_));
  NAND2_X1  g0484(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g0485(.A(new_n525_), .B1(G18), .B2(G178), .ZN(new_n864_));
  INV_X1    g0486(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g0487(.A(G85), .ZN(new_n866_));
  OAI21_X1  g0488(.A(KEYINPUT25), .B1(new_n866_), .B2(G18), .ZN(new_n867_));
  INV_X1    g0489(.A(KEYINPUT25), .ZN(new_n868_));
  NAND3_X1  g0490(.A1(new_n868_), .A2(new_n437_), .A3(G85), .ZN(new_n869_));
  OAI211_X1 g0491(.A(new_n867_), .B(new_n869_), .C1(new_n437_), .C2(G2230), .ZN(new_n870_));
  NAND2_X1  g0492(.A1(new_n865_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g0493(.A(new_n447_), .B1(new_n437_), .B2(G177), .ZN(new_n872_));
  INV_X1    g0494(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g0495(.A1(G18), .A2(G64), .ZN(new_n874_));
  AOI21_X1  g0496(.A(new_n874_), .B1(G18), .B2(G2236), .ZN(new_n875_));
  NAND2_X1  g0497(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g0498(.A1(G18), .A2(G84), .ZN(new_n877_));
  AOI21_X1  g0499(.A(new_n877_), .B1(G18), .B2(G2224), .ZN(new_n878_));
  NAND2_X1  g0500(.A1(G18), .A2(G179), .ZN(new_n879_));
  OAI21_X1  g0501(.A(new_n879_), .B1(new_n529_), .B2(G18), .ZN(new_n880_));
  XNOR2_X1  g0502(.A(new_n878_), .B(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g0503(.A(new_n881_), .B(KEYINPUT26), .ZN(new_n882_));
  NOR2_X1   g0504(.A1(new_n544_), .A2(G18), .ZN(new_n883_));
  AOI21_X1  g0505(.A(new_n883_), .B1(G18), .B2(G180), .ZN(new_n884_));
  NAND2_X1  g0506(.A1(new_n437_), .A2(G83), .ZN(new_n885_));
  OR2_X1    g0507(.A1(new_n885_), .A2(KEYINPUT27), .ZN(new_n886_));
  OAI211_X1 g0508(.A(new_n885_), .B(KEYINPUT27), .C1(new_n437_), .C2(G2218), .ZN(new_n887_));
  NAND2_X1  g0509(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g0510(.A(new_n882_), .B1(new_n884_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g0511(.A(new_n888_), .ZN(new_n890_));
  INV_X1    g0512(.A(new_n884_), .ZN(new_n891_));
  NAND2_X1  g0513(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g0514(.A1(G18), .A2(G65), .ZN(new_n893_));
  AOI21_X1  g0515(.A(new_n893_), .B1(G18), .B2(G2211), .ZN(new_n894_));
  INV_X1    g0516(.A(G171), .ZN(new_n895_));
  OAI21_X1  g0517(.A(new_n555_), .B1(new_n437_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g0518(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g0519(.A1(new_n892_), .A2(new_n897_), .ZN(new_n898_));
  AOI22_X1  g0520(.A1(new_n889_), .A2(new_n898_), .B1(new_n880_), .B2(new_n878_), .ZN(new_n899_));
  NOR2_X1   g0521(.A1(new_n865_), .A2(new_n870_), .ZN(new_n900_));
  OAI211_X1 g0522(.A(new_n871_), .B(new_n876_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n901_));
  AND2_X1   g0523(.A1(new_n856_), .A2(new_n858_), .ZN(new_n902_));
  NOR4_X1   g0524(.A1(new_n852_), .A2(new_n854_), .A3(new_n859_), .A4(new_n902_), .ZN(new_n903_));
  OR2_X1    g0525(.A1(new_n873_), .A2(new_n875_), .ZN(new_n904_));
  AND2_X1   g0526(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g0527(.A(new_n863_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g0528(.A(new_n691_), .ZN(new_n907_));
  AOI21_X1  g0529(.A(new_n907_), .B1(G18), .B2(G189), .ZN(new_n908_));
  NOR2_X1   g0530(.A1(G18), .A2(G62), .ZN(new_n909_));
  AOI21_X1  g0531(.A(new_n909_), .B1(G18), .B2(G4437), .ZN(new_n910_));
  INV_X1    g0532(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g0533(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g0534(.A(new_n684_), .ZN(new_n913_));
  AOI21_X1  g0535(.A(new_n913_), .B1(G18), .B2(G190), .ZN(new_n914_));
  INV_X1    g0536(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g0537(.A1(G18), .A2(G61), .ZN(new_n916_));
  AOI21_X1  g0538(.A(new_n916_), .B1(G18), .B2(G4432), .ZN(new_n917_));
  AND2_X1   g0539(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g0540(.A1(new_n908_), .A2(new_n911_), .ZN(new_n919_));
  AOI21_X1  g0541(.A(new_n912_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g0542(.A(new_n914_), .B(new_n917_), .ZN(new_n921_));
  INV_X1    g0543(.A(new_n656_), .ZN(new_n922_));
  AOI21_X1  g0544(.A(new_n922_), .B1(G18), .B2(G191), .ZN(new_n923_));
  INV_X1    g0545(.A(new_n923_), .ZN(new_n924_));
  NOR2_X1   g0546(.A1(G18), .A2(G60), .ZN(new_n925_));
  AOI21_X1  g0547(.A(new_n925_), .B1(G18), .B2(G4427), .ZN(new_n926_));
  NAND3_X1  g0548(.A1(new_n921_), .A2(new_n924_), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g0549(.A(new_n912_), .ZN(new_n928_));
  NAND2_X1  g0550(.A1(new_n928_), .A2(new_n919_), .ZN(new_n929_));
  OR2_X1    g0551(.A1(new_n924_), .A2(new_n926_), .ZN(new_n930_));
  NAND2_X1  g0552(.A1(new_n924_), .A2(new_n926_), .ZN(new_n931_));
  NAND4_X1  g0553(.A1(new_n930_), .A2(new_n919_), .A3(new_n928_), .A4(new_n931_), .ZN(new_n932_));
  INV_X1    g0554(.A(new_n676_), .ZN(new_n933_));
  AOI21_X1  g0555(.A(new_n933_), .B1(G18), .B2(G192), .ZN(new_n934_));
  INV_X1    g0556(.A(new_n934_), .ZN(new_n935_));
  NOR2_X1   g0557(.A1(G18), .A2(G79), .ZN(new_n936_));
  AOI21_X1  g0558(.A(new_n936_), .B1(G18), .B2(G4420), .ZN(new_n937_));
  NAND3_X1  g0559(.A1(new_n921_), .A2(new_n935_), .A3(new_n937_), .ZN(new_n938_));
  OAI221_X1 g0560(.A(new_n920_), .B1(new_n927_), .B2(new_n929_), .C1(new_n932_), .C2(new_n938_), .ZN(new_n939_));
  INV_X1    g0561(.A(G193), .ZN(new_n940_));
  NOR2_X1   g0562(.A1(new_n940_), .A2(KEYINPUT28), .ZN(new_n941_));
  INV_X1    g0563(.A(new_n941_), .ZN(new_n942_));
  AOI21_X1  g0564(.A(new_n437_), .B1(KEYINPUT28), .B2(new_n940_), .ZN(new_n943_));
  AOI22_X1  g0565(.A1(new_n942_), .A2(new_n943_), .B1(new_n437_), .B2(G47), .ZN(new_n944_));
  NOR2_X1   g0566(.A1(G18), .A2(G80), .ZN(new_n945_));
  AOI21_X1  g0567(.A(new_n945_), .B1(G18), .B2(G4415), .ZN(new_n946_));
  INV_X1    g0568(.A(new_n946_), .ZN(new_n947_));
  NOR2_X1   g0569(.A1(new_n944_), .A2(new_n947_), .ZN(new_n948_));
  INV_X1    g0570(.A(new_n948_), .ZN(new_n949_));
  NAND2_X1  g0571(.A1(new_n944_), .A2(new_n947_), .ZN(new_n950_));
  INV_X1    g0572(.A(new_n950_), .ZN(new_n951_));
  NOR2_X1   g0573(.A1(G18), .A2(G81), .ZN(new_n952_));
  AOI21_X1  g0574(.A(new_n952_), .B1(G18), .B2(G4410), .ZN(new_n953_));
  INV_X1    g0575(.A(G194), .ZN(new_n954_));
  OAI21_X1  g0576(.A(new_n711_), .B1(new_n437_), .B2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g0577(.A1(new_n953_), .A2(new_n955_), .ZN(new_n956_));
  OR2_X1    g0578(.A1(new_n953_), .A2(new_n955_), .ZN(new_n957_));
  NAND4_X1  g0579(.A1(new_n949_), .A2(new_n950_), .A3(new_n956_), .A4(new_n957_), .ZN(new_n958_));
  INV_X1    g0580(.A(G195), .ZN(new_n959_));
  AOI21_X1  g0581(.A(new_n437_), .B1(KEYINPUT29), .B2(new_n959_), .ZN(new_n960_));
  OAI21_X1  g0582(.A(new_n960_), .B1(KEYINPUT29), .B2(new_n959_), .ZN(new_n961_));
  NAND2_X1  g0583(.A1(new_n961_), .A2(new_n721_), .ZN(new_n962_));
  NOR2_X1   g0584(.A1(G18), .A2(G59), .ZN(new_n963_));
  AOI21_X1  g0585(.A(new_n963_), .B1(G18), .B2(G4405), .ZN(new_n964_));
  NAND2_X1  g0586(.A1(new_n962_), .A2(new_n964_), .ZN(new_n965_));
  OAI221_X1 g0587(.A(new_n949_), .B1(new_n951_), .B2(new_n956_), .C1(new_n958_), .C2(new_n965_), .ZN(new_n966_));
  OR2_X1    g0588(.A1(new_n962_), .A2(new_n964_), .ZN(new_n967_));
  INV_X1    g0589(.A(G196), .ZN(new_n968_));
  OAI21_X1  g0590(.A(new_n702_), .B1(new_n437_), .B2(new_n968_), .ZN(new_n969_));
  NAND2_X1  g0591(.A1(new_n700_), .A2(G18), .ZN(new_n970_));
  AOI22_X1  g0592(.A1(new_n970_), .A2(KEYINPUT30), .B1(new_n437_), .B2(G78), .ZN(new_n971_));
  OAI21_X1  g0593(.A(new_n971_), .B1(KEYINPUT30), .B2(new_n970_), .ZN(new_n972_));
  OAI211_X1 g0594(.A(new_n967_), .B(new_n965_), .C1(new_n969_), .C2(new_n972_), .ZN(new_n973_));
  NOR2_X1   g0595(.A1(new_n973_), .A2(new_n958_), .ZN(new_n974_));
  NAND2_X1  g0596(.A1(new_n972_), .A2(new_n969_), .ZN(new_n975_));
  NOR2_X1   g0597(.A1(G18), .A2(G77), .ZN(new_n976_));
  AOI21_X1  g0598(.A(new_n976_), .B1(G18), .B2(G4394), .ZN(new_n977_));
  INV_X1    g0599(.A(G187), .ZN(new_n978_));
  OAI21_X1  g0600(.A(new_n705_), .B1(new_n437_), .B2(new_n978_), .ZN(new_n979_));
  NAND2_X1  g0601(.A1(new_n977_), .A2(new_n979_), .ZN(new_n980_));
  AND2_X1   g0602(.A1(new_n975_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1    g0603(.A(new_n981_), .ZN(new_n982_));
  AOI21_X1  g0604(.A(new_n966_), .B1(new_n974_), .B2(new_n982_), .ZN(new_n983_));
  INV_X1    g0605(.A(new_n592_), .ZN(new_n984_));
  AOI21_X1  g0606(.A(new_n984_), .B1(G18), .B2(G203), .ZN(new_n985_));
  INV_X1    g0607(.A(new_n985_), .ZN(new_n986_));
  NOR2_X1   g0608(.A1(G18), .A2(G53), .ZN(new_n987_));
  AOI21_X1  g0609(.A(new_n987_), .B1(G18), .B2(G3729), .ZN(new_n988_));
  INV_X1    g0610(.A(G202), .ZN(new_n989_));
  OAI21_X1  g0611(.A(new_n601_), .B1(new_n437_), .B2(new_n989_), .ZN(new_n990_));
  NOR2_X1   g0612(.A1(G18), .A2(G54), .ZN(new_n991_));
  AOI21_X1  g0613(.A(new_n991_), .B1(G18), .B2(G3737), .ZN(new_n992_));
  AOI22_X1  g0614(.A1(new_n986_), .A2(new_n988_), .B1(new_n990_), .B2(new_n992_), .ZN(new_n993_));
  OAI21_X1  g0615(.A(new_n993_), .B1(new_n986_), .B2(new_n988_), .ZN(new_n994_));
  NOR2_X1   g0616(.A1(G18), .A2(G55), .ZN(new_n995_));
  AOI21_X1  g0617(.A(new_n995_), .B1(G18), .B2(G3743), .ZN(new_n996_));
  INV_X1    g0618(.A(G201), .ZN(new_n997_));
  OAI21_X1  g0619(.A(new_n608_), .B1(new_n437_), .B2(new_n997_), .ZN(new_n998_));
  NAND2_X1  g0620(.A1(new_n996_), .A2(new_n998_), .ZN(new_n999_));
  AOI21_X1  g0621(.A(new_n614_), .B1(G18), .B2(G200), .ZN(new_n1000_));
  NAND2_X1  g0622(.A1(G18), .A2(G3749), .ZN(new_n1001_));
  OAI21_X1  g0623(.A(new_n1001_), .B1(G18), .B2(G56), .ZN(new_n1002_));
  OAI21_X1  g0624(.A(new_n999_), .B1(new_n1000_), .B2(new_n1002_), .ZN(new_n1003_));
  NAND2_X1  g0625(.A1(new_n1000_), .A2(new_n1002_), .ZN(new_n1004_));
  OAI221_X1 g0626(.A(new_n1004_), .B1(new_n998_), .B2(new_n996_), .C1(new_n990_), .C2(new_n992_), .ZN(new_n1005_));
  NOR3_X1   g0627(.A1(new_n994_), .A2(new_n1003_), .A3(new_n1005_), .ZN(new_n1006_));
  MUX2_X1   g0628(.A(G103), .B(G204), .S(G18), .Z(new_n1007_));
  NOR2_X1   g0629(.A1(G18), .A2(G73), .ZN(new_n1008_));
  AOI21_X1  g0630(.A(new_n1008_), .B1(G18), .B2(G3723), .ZN(new_n1009_));
  OR2_X1    g0631(.A1(new_n1007_), .A2(new_n1009_), .ZN(new_n1010_));
  INV_X1    g0632(.A(new_n1010_), .ZN(new_n1011_));
  AND2_X1   g0633(.A1(new_n437_), .A2(G75), .ZN(new_n1012_));
  NOR2_X1   g0634(.A1(new_n437_), .A2(G3717), .ZN(new_n1013_));
  OAI21_X1  g0635(.A(KEYINPUT20), .B1(new_n1012_), .B2(new_n1013_), .ZN(new_n1014_));
  OAI21_X1  g0636(.A(new_n1014_), .B1(KEYINPUT20), .B2(new_n1013_), .ZN(new_n1015_));
  NOR2_X1   g0637(.A1(new_n638_), .A2(G18), .ZN(new_n1016_));
  AOI21_X1  g0638(.A(new_n1016_), .B1(G18), .B2(G205), .ZN(new_n1017_));
  INV_X1    g0639(.A(new_n1017_), .ZN(new_n1018_));
  NOR2_X1   g0640(.A1(new_n1015_), .A2(new_n1018_), .ZN(new_n1019_));
  INV_X1    g0641(.A(G206), .ZN(new_n1020_));
  OAI21_X1  g0642(.A(new_n753_), .B1(new_n437_), .B2(new_n1020_), .ZN(new_n1021_));
  XNOR2_X1  g0643(.A(new_n1021_), .B(KEYINPUT21), .ZN(new_n1022_));
  NOR2_X1   g0644(.A1(G18), .A2(G76), .ZN(new_n1023_));
  AOI21_X1  g0645(.A(new_n1023_), .B1(G18), .B2(G3711), .ZN(new_n1024_));
  INV_X1    g0646(.A(new_n1024_), .ZN(new_n1025_));
  AOI21_X1  g0647(.A(new_n1019_), .B1(new_n1022_), .B2(new_n1025_), .ZN(new_n1026_));
  NOR2_X1   g0648(.A1(G18), .A2(G74), .ZN(new_n1027_));
  AOI21_X1  g0649(.A(new_n1027_), .B1(G18), .B2(G3705), .ZN(new_n1028_));
  INV_X1    g0650(.A(G207), .ZN(new_n1029_));
  OAI21_X1  g0651(.A(new_n758_), .B1(new_n437_), .B2(new_n1029_), .ZN(new_n1030_));
  NAND2_X1  g0652(.A1(new_n1028_), .A2(new_n1030_), .ZN(new_n1031_));
  NOR2_X1   g0653(.A1(new_n1028_), .A2(new_n1030_), .ZN(new_n1032_));
  NAND3_X1  g0654(.A1(new_n437_), .A2(G41), .A3(G70), .ZN(new_n1033_));
  OAI21_X1  g0655(.A(new_n1031_), .B1(new_n1032_), .B2(new_n1033_), .ZN(new_n1034_));
  NOR2_X1   g0656(.A1(new_n1022_), .A2(new_n1025_), .ZN(new_n1035_));
  OAI21_X1  g0657(.A(new_n1026_), .B1(new_n1034_), .B2(new_n1035_), .ZN(new_n1036_));
  NAND2_X1  g0658(.A1(new_n1015_), .A2(new_n1018_), .ZN(new_n1037_));
  AOI21_X1  g0659(.A(new_n1011_), .B1(new_n1036_), .B2(new_n1037_), .ZN(new_n1038_));
  AOI21_X1  g0660(.A(new_n1035_), .B1(new_n1018_), .B2(new_n1015_), .ZN(new_n1039_));
  INV_X1    g0661(.A(new_n1032_), .ZN(new_n1040_));
  NAND2_X1  g0662(.A1(new_n1007_), .A2(new_n1009_), .ZN(new_n1041_));
  NAND4_X1  g0663(.A1(new_n1040_), .A2(new_n1010_), .A3(new_n1031_), .A4(new_n1041_), .ZN(new_n1042_));
  NAND2_X1  g0664(.A1(new_n437_), .A2(G41), .ZN(new_n1043_));
  NOR2_X1   g0665(.A1(G18), .A2(G70), .ZN(new_n1044_));
  NAND2_X1  g0666(.A1(new_n1043_), .A2(new_n1044_), .ZN(new_n1045_));
  NAND3_X1  g0667(.A1(new_n1045_), .A2(G89), .A3(new_n1033_), .ZN(new_n1046_));
  NOR2_X1   g0668(.A1(new_n1042_), .A2(new_n1046_), .ZN(new_n1047_));
  NAND3_X1  g0669(.A1(new_n1039_), .A2(new_n1026_), .A3(new_n1047_), .ZN(new_n1048_));
  NAND2_X1  g0670(.A1(new_n1048_), .A2(new_n1041_), .ZN(new_n1049_));
  OAI21_X1  g0671(.A(new_n1006_), .B1(new_n1038_), .B2(new_n1049_), .ZN(new_n1050_));
  NOR3_X1   g0672(.A1(new_n1005_), .A2(new_n1003_), .A3(new_n993_), .ZN(new_n1051_));
  AOI21_X1  g0673(.A(new_n1051_), .B1(new_n1003_), .B2(new_n1004_), .ZN(new_n1052_));
  AND2_X1   g0674(.A1(new_n1050_), .A2(new_n1052_), .ZN(new_n1053_));
  OAI211_X1 g0675(.A(new_n974_), .B(new_n981_), .C1(new_n979_), .C2(new_n977_), .ZN(new_n1054_));
  OAI21_X1  g0676(.A(new_n983_), .B1(new_n1053_), .B2(new_n1054_), .ZN(new_n1055_));
  OR2_X1    g0677(.A1(new_n935_), .A2(new_n937_), .ZN(new_n1056_));
  NAND2_X1  g0678(.A1(new_n935_), .A2(new_n937_), .ZN(new_n1057_));
  NAND3_X1  g0679(.A1(new_n921_), .A2(new_n1056_), .A3(new_n1057_), .ZN(new_n1058_));
  NOR2_X1   g0680(.A1(new_n932_), .A2(new_n1058_), .ZN(new_n1059_));
  AOI21_X1  g0681(.A(new_n939_), .B1(new_n1055_), .B2(new_n1059_), .ZN(new_n1060_));
  INV_X1    g0682(.A(new_n892_), .ZN(new_n1061_));
  OR2_X1    g0683(.A1(new_n894_), .A2(new_n896_), .ZN(new_n1062_));
  NAND4_X1  g0684(.A1(new_n904_), .A2(new_n1062_), .A3(new_n876_), .A4(new_n897_), .ZN(new_n1063_));
  INV_X1    g0685(.A(new_n871_), .ZN(new_n1064_));
  NOR4_X1   g0686(.A1(new_n1061_), .A2(new_n1063_), .A3(new_n1064_), .A4(new_n900_), .ZN(new_n1065_));
  NAND3_X1  g0687(.A1(new_n889_), .A2(new_n903_), .A3(new_n1065_), .ZN(new_n1066_));
  OAI21_X1  g0688(.A(new_n906_), .B1(new_n1060_), .B2(new_n1066_), .ZN(new_n1067_));
  AOI21_X1  g0689(.A(new_n820_), .B1(new_n511_), .B2(new_n822_), .ZN(new_n1068_));
  NOR2_X1   g0690(.A1(new_n813_), .A2(new_n819_), .ZN(new_n1069_));
  NAND3_X1  g0691(.A1(new_n1068_), .A2(new_n1069_), .A3(new_n830_), .ZN(new_n1070_));
  NOR3_X1   g0692(.A1(new_n1070_), .A2(new_n808_), .A3(new_n828_), .ZN(new_n1071_));
  AOI21_X1  g0693(.A(new_n832_), .B1(new_n1067_), .B2(new_n1071_), .ZN(new_n1072_));
  NAND2_X1  g0694(.A1(new_n801_), .A2(G38), .ZN(new_n1073_));
  XNOR2_X1  g0695(.A(new_n802_), .B(KEYINPUT23), .ZN(new_n1074_));
  AND2_X1   g0696(.A1(new_n1074_), .A2(new_n801_), .ZN(new_n1075_));
  INV_X1    g0697(.A(G38), .ZN(new_n1076_));
  NOR2_X1   g0698(.A1(new_n1074_), .A2(new_n1076_), .ZN(new_n1077_));
  OAI21_X1  g0699(.A(new_n1073_), .B1(new_n1075_), .B2(new_n1077_), .ZN(new_n1078_));
  OAI21_X1  g0700(.A(new_n803_), .B1(new_n1072_), .B2(new_n1078_), .ZN(G258));
  OAI21_X1  g0701(.A(new_n803_), .B1(new_n1072_), .B2(new_n1078_), .ZN(G264));
  NAND4_X1  g0702(.A1(new_n769_), .A2(new_n775_), .A3(new_n732_), .A4(new_n795_), .ZN(new_n1081_));
  NOR2_X1   g0703(.A1(new_n581_), .A2(new_n589_), .ZN(new_n1082_));
  AOI21_X1  g0704(.A(new_n582_), .B1(new_n1081_), .B2(new_n1082_), .ZN(new_n1083_));
  XOR2_X1   g0705(.A(new_n459_), .B(KEYINPUT31), .Z(new_n1084_));
  NAND2_X1  g0706(.A1(new_n1084_), .A2(new_n741_), .ZN(new_n1085_));
  NAND2_X1  g0707(.A1(new_n737_), .A2(new_n739_), .ZN(new_n1086_));
  NOR3_X1   g0708(.A1(new_n1085_), .A2(new_n1086_), .A3(new_n466_), .ZN(new_n1087_));
  XNOR2_X1  g0709(.A(new_n1087_), .B(KEYINPUT32), .ZN(new_n1088_));
  INV_X1    g0710(.A(new_n1088_), .ZN(new_n1089_));
  OAI21_X1  g0711(.A(new_n487_), .B1(new_n1083_), .B2(new_n1089_), .ZN(new_n1090_));
  INV_X1    g0712(.A(new_n1090_), .ZN(new_n1091_));
  OAI21_X1  g0713(.A(new_n446_), .B1(new_n1091_), .B2(new_n494_), .ZN(G270));
  INV_X1    g0714(.A(new_n766_), .ZN(new_n1093_));
  INV_X1    g0715(.A(new_n644_), .ZN(new_n1094_));
  NAND2_X1  g0716(.A1(new_n652_), .A2(G4526), .ZN(new_n1095_));
  OAI21_X1  g0717(.A(new_n1093_), .B1(new_n1094_), .B2(new_n1095_), .ZN(new_n1096_));
  XNOR2_X1  g0718(.A(new_n1096_), .B(new_n628_), .ZN(G388));
  NAND2_X1  g0719(.A1(new_n756_), .A2(new_n755_), .ZN(new_n1098_));
  AOI21_X1  g0720(.A(new_n761_), .B1(new_n759_), .B2(new_n1098_), .ZN(new_n1099_));
  NAND3_X1  g0721(.A1(new_n649_), .A2(new_n762_), .A3(new_n650_), .ZN(new_n1100_));
  OAI21_X1  g0722(.A(new_n1099_), .B1(new_n636_), .B2(new_n1100_), .ZN(new_n1101_));
  INV_X1    g0723(.A(G4526), .ZN(new_n1102_));
  NOR2_X1   g0724(.A1(new_n439_), .A2(new_n1102_), .ZN(new_n1103_));
  NOR2_X1   g0725(.A1(new_n636_), .A2(new_n651_), .ZN(new_n1104_));
  AOI21_X1  g0726(.A(new_n1101_), .B1(new_n1103_), .B2(new_n1104_), .ZN(new_n1105_));
  XNOR2_X1  g0727(.A(new_n1105_), .B(new_n752_), .ZN(G391));
  NAND2_X1  g0728(.A1(new_n1100_), .A2(new_n649_), .ZN(new_n1107_));
  INV_X1    g0729(.A(new_n1107_), .ZN(new_n1108_));
  NAND2_X1  g0730(.A1(new_n1095_), .A2(new_n1108_), .ZN(new_n1109_));
  NOR2_X1   g0731(.A1(new_n635_), .A2(new_n632_), .ZN(new_n1110_));
  NOR2_X1   g0732(.A1(new_n761_), .A2(new_n1110_), .ZN(new_n1111_));
  INV_X1    g0733(.A(new_n1111_), .ZN(new_n1112_));
  XNOR2_X1  g0734(.A(new_n1109_), .B(new_n1112_), .ZN(G394));
  NOR2_X1   g0735(.A1(new_n1103_), .A2(new_n762_), .ZN(new_n1114_));
  INV_X1    g0736(.A(new_n651_), .ZN(new_n1115_));
  XNOR2_X1  g0737(.A(new_n1114_), .B(new_n1115_), .ZN(G397));
  NAND2_X1  g0738(.A1(new_n767_), .A2(new_n653_), .ZN(new_n1117_));
  NAND2_X1  g0739(.A1(new_n596_), .A2(new_n605_), .ZN(new_n1118_));
  NAND3_X1  g0740(.A1(new_n611_), .A2(new_n1118_), .A3(new_n748_), .ZN(new_n1119_));
  AND2_X1   g0741(.A1(new_n1119_), .A2(new_n612_), .ZN(new_n1120_));
  INV_X1    g0742(.A(new_n1120_), .ZN(new_n1121_));
  NAND2_X1  g0743(.A1(new_n1117_), .A2(new_n1121_), .ZN(new_n1122_));
  INV_X1    g0744(.A(new_n749_), .ZN(new_n1123_));
  NAND2_X1  g0745(.A1(new_n1123_), .A2(new_n611_), .ZN(new_n1124_));
  AND2_X1   g0746(.A1(new_n1124_), .A2(new_n612_), .ZN(new_n1125_));
  OAI21_X1  g0747(.A(new_n1122_), .B1(new_n1117_), .B2(new_n1125_), .ZN(new_n1126_));
  XOR2_X1   g0748(.A(new_n1126_), .B(new_n618_), .Z(G376));
  AOI21_X1  g0749(.A(new_n749_), .B1(new_n1117_), .B2(new_n607_), .ZN(new_n1128_));
  XOR2_X1   g0750(.A(new_n1128_), .B(new_n613_), .Z(G379));
  INV_X1    g0751(.A(new_n1117_), .ZN(new_n1130_));
  NAND2_X1  g0752(.A1(new_n1130_), .A2(new_n747_), .ZN(new_n1131_));
  OAI21_X1  g0753(.A(new_n1131_), .B1(new_n596_), .B2(new_n1130_), .ZN(new_n1132_));
  NOR2_X1   g0754(.A1(new_n606_), .A2(new_n604_), .ZN(new_n1133_));
  XNOR2_X1  g0755(.A(new_n1132_), .B(new_n1133_), .ZN(G382));
  XNOR2_X1  g0756(.A(new_n1117_), .B(new_n600_), .ZN(G385));
  INV_X1    g0757(.A(G229), .ZN(new_n1136_));
  OAI21_X1  g0758(.A(new_n1043_), .B1(new_n437_), .B2(new_n1136_), .ZN(new_n1137_));
  XNOR2_X1  g0759(.A(new_n1137_), .B(new_n632_), .ZN(new_n1138_));
  XNOR2_X1  g0760(.A(new_n1138_), .B(new_n647_), .ZN(new_n1139_));
  NAND2_X1  g0761(.A1(new_n437_), .A2(G44), .ZN(new_n1140_));
  INV_X1    g0762(.A(new_n1140_), .ZN(new_n1141_));
  AOI21_X1  g0763(.A(new_n1141_), .B1(G18), .B2(G239), .ZN(new_n1142_));
  AOI21_X1  g0764(.A(KEYINPUT33), .B1(new_n1139_), .B2(new_n1142_), .ZN(new_n1143_));
  OAI21_X1  g0765(.A(new_n1143_), .B1(new_n1142_), .B2(new_n1139_), .ZN(new_n1144_));
  XNOR2_X1  g0766(.A(new_n1144_), .B(new_n625_), .ZN(new_n1145_));
  XNOR2_X1  g0767(.A(new_n610_), .B(new_n595_), .ZN(new_n1146_));
  XNOR2_X1  g0768(.A(new_n615_), .B(new_n603_), .ZN(new_n1147_));
  XNOR2_X1  g0769(.A(new_n1146_), .B(new_n1147_), .ZN(new_n1148_));
  XNOR2_X1  g0770(.A(new_n1148_), .B(new_n639_), .ZN(new_n1149_));
  XNOR2_X1  g0771(.A(new_n1145_), .B(new_n1149_), .ZN(new_n1150_));
  NAND2_X1  g0772(.A1(new_n447_), .A2(G18), .ZN(new_n1151_));
  INV_X1    g0773(.A(G211), .ZN(new_n1152_));
  OR2_X1    g0774(.A1(new_n1152_), .A2(G212), .ZN(new_n1153_));
  NAND2_X1  g0775(.A1(new_n1152_), .A2(G212), .ZN(new_n1154_));
  AOI21_X1  g0776(.A(new_n1151_), .B1(new_n1153_), .B2(new_n1154_), .ZN(new_n1155_));
  NOR2_X1   g0777(.A1(new_n1155_), .A2(new_n511_), .ZN(new_n1156_));
  XOR2_X1   g0778(.A(new_n454_), .B(new_n475_), .Z(new_n1157_));
  XNOR2_X1  g0779(.A(new_n1157_), .B(new_n469_), .ZN(new_n1158_));
  NOR2_X1   g0780(.A1(new_n437_), .A2(G215), .ZN(new_n1159_));
  XOR2_X1   g0781(.A(new_n462_), .B(new_n1159_), .Z(new_n1160_));
  XNOR2_X1  g0782(.A(new_n1158_), .B(new_n1160_), .ZN(new_n1161_));
  MUX2_X1   g0783(.A(new_n1155_), .B(new_n1156_), .S(new_n1161_), .Z(new_n1162_));
  XNOR2_X1  g0784(.A(new_n557_), .B(new_n545_), .ZN(new_n1163_));
  INV_X1    g0785(.A(G141), .ZN(new_n1164_));
  NOR2_X1   g0786(.A1(new_n1164_), .A2(G18), .ZN(new_n1165_));
  AOI21_X1  g0787(.A(new_n1165_), .B1(G18), .B2(G161), .ZN(new_n1166_));
  XNOR2_X1  g0788(.A(new_n1163_), .B(new_n1166_), .ZN(new_n1167_));
  XNOR2_X1  g0789(.A(new_n566_), .B(new_n526_), .ZN(new_n1168_));
  XNOR2_X1  g0790(.A(new_n1167_), .B(new_n1168_), .ZN(new_n1169_));
  XOR2_X1   g0791(.A(new_n502_), .B(new_n533_), .Z(new_n1170_));
  XNOR2_X1  g0792(.A(new_n1169_), .B(new_n1170_), .ZN(new_n1171_));
  NAND3_X1  g0793(.A1(new_n506_), .A2(G18), .A3(new_n512_), .ZN(new_n1172_));
  INV_X1    g0794(.A(new_n513_), .ZN(new_n1173_));
  OAI21_X1  g0795(.A(new_n1172_), .B1(new_n1173_), .B2(new_n505_), .ZN(new_n1174_));
  XOR2_X1   g0796(.A(new_n1174_), .B(new_n497_), .Z(new_n1175_));
  AOI21_X1  g0797(.A(new_n1162_), .B1(new_n1171_), .B2(new_n1175_), .ZN(new_n1176_));
  OAI21_X1  g0798(.A(new_n1176_), .B1(new_n1175_), .B2(new_n1171_), .ZN(new_n1177_));
  XOR2_X1   g0799(.A(new_n725_), .B(new_n778_), .Z(new_n1178_));
  XOR2_X1   g0800(.A(new_n699_), .B(new_n786_), .Z(new_n1179_));
  OR2_X1    g0801(.A1(new_n1178_), .A2(new_n1179_), .ZN(new_n1180_));
  NAND2_X1  g0802(.A1(new_n437_), .A2(G115), .ZN(new_n1181_));
  INV_X1    g0803(.A(G227), .ZN(new_n1182_));
  OAI21_X1  g0804(.A(new_n1181_), .B1(new_n437_), .B2(new_n1182_), .ZN(new_n1183_));
  INV_X1    g0805(.A(G118), .ZN(new_n1184_));
  OAI21_X1  g0806(.A(new_n706_), .B1(new_n1184_), .B2(G18), .ZN(new_n1185_));
  XNOR2_X1  g0807(.A(new_n1183_), .B(new_n1185_), .ZN(new_n1186_));
  NOR2_X1   g0808(.A1(new_n1180_), .A2(new_n1186_), .ZN(new_n1187_));
  XOR2_X1   g0809(.A(new_n1187_), .B(KEYINPUT35), .Z(new_n1188_));
  NAND2_X1  g0810(.A1(new_n1178_), .A2(new_n1179_), .ZN(new_n1189_));
  NOR2_X1   g0811(.A1(new_n1189_), .A2(new_n1186_), .ZN(new_n1190_));
  XNOR2_X1  g0812(.A(new_n1190_), .B(KEYINPUT34), .ZN(new_n1191_));
  NAND3_X1  g0813(.A1(new_n1180_), .A2(new_n1186_), .A3(new_n1189_), .ZN(new_n1192_));
  NAND3_X1  g0814(.A1(new_n1188_), .A2(new_n1191_), .A3(new_n1192_), .ZN(new_n1193_));
  XNOR2_X1  g0815(.A(new_n1193_), .B(new_n687_), .ZN(new_n1194_));
  XNOR2_X1  g0816(.A(new_n1194_), .B(new_n662_), .ZN(new_n1195_));
  XNOR2_X1  g0817(.A(new_n693_), .B(new_n678_), .ZN(new_n1196_));
  AOI211_X1 g0818(.A(new_n1150_), .B(new_n1177_), .C1(new_n1195_), .C2(new_n1196_), .ZN(new_n1197_));
  OR2_X1    g0819(.A1(new_n1195_), .A2(new_n1196_), .ZN(new_n1198_));
  NAND2_X1  g0820(.A1(new_n1197_), .A2(new_n1198_), .ZN(G412));
  XOR2_X1   g0821(.A(new_n1009_), .B(new_n1028_), .Z(new_n1200_));
  XNOR2_X1  g0822(.A(new_n1200_), .B(new_n1015_), .ZN(new_n1201_));
  NAND2_X1  g0823(.A1(new_n437_), .A2(G69), .ZN(new_n1202_));
  OAI21_X1  g0824(.A(new_n1202_), .B1(new_n437_), .B2(G3698), .ZN(new_n1203_));
  XNOR2_X1  g0825(.A(new_n1201_), .B(new_n1203_), .ZN(new_n1204_));
  AOI21_X1  g0826(.A(new_n1044_), .B1(G18), .B2(G3701), .ZN(new_n1205_));
  XNOR2_X1  g0827(.A(new_n1024_), .B(new_n1205_), .ZN(new_n1206_));
  XNOR2_X1  g0828(.A(new_n1204_), .B(new_n1206_), .ZN(new_n1207_));
  XNOR2_X1  g0829(.A(new_n992_), .B(new_n1002_), .ZN(new_n1208_));
  XNOR2_X1  g0830(.A(new_n1207_), .B(new_n1208_), .ZN(new_n1209_));
  XOR2_X1   g0831(.A(new_n996_), .B(new_n988_), .Z(new_n1210_));
  XNOR2_X1  g0832(.A(new_n1209_), .B(new_n1210_), .ZN(new_n1211_));
  XOR2_X1   g0833(.A(new_n964_), .B(new_n977_), .Z(new_n1212_));
  XNOR2_X1  g0834(.A(new_n1212_), .B(new_n972_), .ZN(new_n1213_));
  XNOR2_X1  g0835(.A(new_n1213_), .B(new_n947_), .ZN(new_n1214_));
  XNOR2_X1  g0836(.A(new_n910_), .B(new_n926_), .ZN(new_n1215_));
  XNOR2_X1  g0837(.A(new_n1215_), .B(new_n917_), .ZN(new_n1216_));
  XNOR2_X1  g0838(.A(new_n1214_), .B(new_n1216_), .ZN(new_n1217_));
  NAND2_X1  g0839(.A1(G18), .A2(G4393), .ZN(new_n1218_));
  OAI21_X1  g0840(.A(new_n1218_), .B1(G18), .B2(G58), .ZN(new_n1219_));
  XNOR2_X1  g0841(.A(new_n953_), .B(new_n1219_), .ZN(new_n1220_));
  XNOR2_X1  g0842(.A(new_n1220_), .B(new_n937_), .ZN(new_n1221_));
  XNOR2_X1  g0843(.A(new_n1217_), .B(new_n1221_), .ZN(new_n1222_));
  XOR2_X1   g0844(.A(new_n878_), .B(new_n875_), .Z(new_n1223_));
  XNOR2_X1  g0845(.A(new_n1223_), .B(new_n870_), .ZN(new_n1224_));
  NAND2_X1  g0846(.A1(new_n437_), .A2(G82), .ZN(new_n1225_));
  OAI21_X1  g0847(.A(new_n1225_), .B1(new_n437_), .B2(G2208), .ZN(new_n1226_));
  XNOR2_X1  g0848(.A(new_n1224_), .B(new_n1226_), .ZN(new_n1227_));
  XNOR2_X1  g0849(.A(new_n840_), .B(new_n847_), .ZN(new_n1228_));
  XOR2_X1   g0850(.A(new_n1228_), .B(new_n858_), .Z(new_n1229_));
  XNOR2_X1  g0851(.A(new_n1227_), .B(new_n1229_), .ZN(new_n1230_));
  XNOR2_X1  g0852(.A(new_n888_), .B(new_n894_), .ZN(new_n1231_));
  XNOR2_X1  g0853(.A(new_n1231_), .B(new_n853_), .ZN(new_n1232_));
  AND2_X1   g0854(.A1(new_n1230_), .A2(new_n1232_), .ZN(new_n1233_));
  NOR2_X1   g0855(.A1(new_n1230_), .A2(new_n1232_), .ZN(new_n1234_));
  XNOR2_X1  g0856(.A(new_n806_), .B(new_n818_), .ZN(new_n1235_));
  XNOR2_X1  g0857(.A(new_n1235_), .B(new_n810_), .ZN(new_n1236_));
  NOR2_X1   g0858(.A1(new_n437_), .A2(G1459), .ZN(new_n1237_));
  AOI21_X1  g0859(.A(new_n1237_), .B1(new_n437_), .B2(G114), .ZN(new_n1238_));
  XNOR2_X1  g0860(.A(new_n1236_), .B(new_n1238_), .ZN(new_n1239_));
  OAI21_X1  g0861(.A(new_n437_), .B1(G1455), .B2(G2204), .ZN(new_n1240_));
  AOI21_X1  g0862(.A(new_n1240_), .B1(G1455), .B2(G2204), .ZN(new_n1241_));
  XOR2_X1   g0863(.A(G1492), .B(G1496), .Z(new_n1242_));
  AOI21_X1  g0864(.A(new_n1241_), .B1(G18), .B2(new_n1242_), .ZN(new_n1243_));
  XNOR2_X1  g0865(.A(new_n822_), .B(new_n824_), .ZN(new_n1244_));
  XNOR2_X1  g0866(.A(new_n1243_), .B(new_n1244_), .ZN(new_n1245_));
  XOR2_X1   g0867(.A(new_n1239_), .B(new_n1245_), .Z(new_n1246_));
  NOR3_X1   g0868(.A1(new_n1233_), .A2(new_n1234_), .A3(new_n1246_), .ZN(new_n1247_));
  NAND3_X1  g0869(.A1(new_n1211_), .A2(new_n1222_), .A3(new_n1247_), .ZN(G414));
  XNOR2_X1  g0870(.A(new_n896_), .B(new_n872_), .ZN(new_n1249_));
  XNOR2_X1  g0871(.A(new_n1249_), .B(new_n865_), .ZN(new_n1250_));
  XNOR2_X1  g0872(.A(new_n1250_), .B(new_n880_), .ZN(new_n1251_));
  OAI21_X1  g0873(.A(G18), .B1(KEYINPUT36), .B2(G181), .ZN(new_n1252_));
  AND2_X1   g0874(.A1(KEYINPUT36), .A2(G181), .ZN(new_n1253_));
  OAI22_X1  g0875(.A1(new_n1252_), .A2(new_n1253_), .B1(G18), .B2(new_n1164_), .ZN(new_n1254_));
  XOR2_X1   g0876(.A(new_n884_), .B(new_n1254_), .Z(new_n1255_));
  MUX2_X1   g0877(.A(new_n841_), .B(new_n850_), .S(new_n856_), .Z(new_n1256_));
  XOR2_X1   g0878(.A(new_n1255_), .B(new_n1256_), .Z(new_n1257_));
  XNOR2_X1  g0879(.A(new_n1251_), .B(new_n1257_), .ZN(new_n1258_));
  NOR2_X1   g0880(.A1(new_n833_), .A2(new_n843_), .ZN(new_n1259_));
  AOI21_X1  g0881(.A(new_n1259_), .B1(new_n845_), .B2(new_n833_), .ZN(new_n1260_));
  INV_X1    g0882(.A(new_n1260_), .ZN(new_n1261_));
  NOR2_X1   g0883(.A1(new_n1258_), .A2(new_n1261_), .ZN(new_n1262_));
  AND2_X1   g0884(.A1(new_n1258_), .A2(new_n1261_), .ZN(new_n1263_));
  XNOR2_X1  g0885(.A(new_n1000_), .B(new_n990_), .ZN(new_n1264_));
  XNOR2_X1  g0886(.A(new_n1264_), .B(new_n986_), .ZN(new_n1265_));
  INV_X1    g0887(.A(G198), .ZN(new_n1266_));
  OAI21_X1  g0888(.A(new_n1043_), .B1(new_n437_), .B2(new_n1266_), .ZN(new_n1267_));
  XOR2_X1   g0889(.A(new_n1007_), .B(new_n1267_), .Z(new_n1268_));
  AOI21_X1  g0890(.A(new_n1141_), .B1(G18), .B2(G208), .ZN(new_n1269_));
  XNOR2_X1  g0891(.A(new_n1268_), .B(new_n1269_), .ZN(new_n1270_));
  XNOR2_X1  g0892(.A(new_n1270_), .B(new_n1030_), .ZN(new_n1271_));
  XNOR2_X1  g0893(.A(new_n1022_), .B(new_n1018_), .ZN(new_n1272_));
  XNOR2_X1  g0894(.A(new_n1272_), .B(new_n998_), .ZN(new_n1273_));
  XNOR2_X1  g0895(.A(new_n1271_), .B(new_n1273_), .ZN(new_n1274_));
  AOI211_X1 g0896(.A(new_n1262_), .B(new_n1263_), .C1(new_n1265_), .C2(new_n1274_), .ZN(new_n1275_));
  INV_X1    g0897(.A(G166), .ZN(new_n1276_));
  AOI21_X1  g0898(.A(new_n812_), .B1(G18), .B2(new_n1276_), .ZN(new_n1277_));
  AOI21_X1  g0899(.A(new_n1277_), .B1(new_n804_), .B2(new_n812_), .ZN(new_n1278_));
  MUX2_X1   g0900(.A(new_n815_), .B(new_n816_), .S(new_n829_), .Z(new_n1279_));
  OR2_X1    g0901(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1280_));
  NAND2_X1  g0902(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1281_));
  NAND3_X1  g0903(.A1(new_n1280_), .A2(KEYINPUT37), .A3(new_n1281_), .ZN(new_n1282_));
  NOR2_X1   g0904(.A1(new_n1151_), .A2(G170), .ZN(new_n1283_));
  XNOR2_X1  g0905(.A(new_n1282_), .B(new_n1283_), .ZN(new_n1284_));
  INV_X1    g0906(.A(G164), .ZN(new_n1285_));
  OR2_X1    g0907(.A1(new_n1285_), .A2(G165), .ZN(new_n1286_));
  NAND2_X1  g0908(.A1(new_n1285_), .A2(G165), .ZN(new_n1287_));
  AOI21_X1  g0909(.A(new_n1151_), .B1(new_n1286_), .B2(new_n1287_), .ZN(new_n1288_));
  XNOR2_X1  g0910(.A(new_n1284_), .B(new_n1288_), .ZN(new_n1289_));
  XNOR2_X1  g0911(.A(new_n944_), .B(new_n969_), .ZN(new_n1290_));
  XNOR2_X1  g0912(.A(new_n1290_), .B(new_n915_), .ZN(new_n1291_));
  XNOR2_X1  g0913(.A(new_n955_), .B(new_n979_), .ZN(new_n1292_));
  INV_X1    g0914(.A(G197), .ZN(new_n1293_));
  OAI21_X1  g0915(.A(new_n1181_), .B1(new_n437_), .B2(new_n1293_), .ZN(new_n1294_));
  XNOR2_X1  g0916(.A(new_n1292_), .B(new_n1294_), .ZN(new_n1295_));
  XNOR2_X1  g0917(.A(new_n1295_), .B(new_n962_), .ZN(new_n1296_));
  XNOR2_X1  g0918(.A(new_n908_), .B(new_n923_), .ZN(new_n1297_));
  XNOR2_X1  g0919(.A(new_n1297_), .B(new_n934_), .ZN(new_n1298_));
  XNOR2_X1  g0920(.A(new_n1296_), .B(new_n1298_), .ZN(new_n1299_));
  AOI21_X1  g0921(.A(new_n1289_), .B1(new_n1291_), .B2(new_n1299_), .ZN(new_n1300_));
  OR2_X1    g0922(.A1(new_n1299_), .A2(new_n1291_), .ZN(new_n1301_));
  OR2_X1    g0923(.A1(new_n1274_), .A2(new_n1265_), .ZN(new_n1302_));
  NAND4_X1  g0924(.A1(new_n1275_), .A2(new_n1300_), .A3(new_n1301_), .A4(new_n1302_), .ZN(G416));
  XNOR2_X1  g0925(.A(G258), .B(KEYINPUT38), .ZN(G249));
  NAND2_X1  g0926(.A1(new_n559_), .A2(new_n584_), .ZN(new_n1305_));
  XNOR2_X1  g0927(.A(new_n1081_), .B(new_n1305_), .ZN(G295));
  NOR2_X1   g0928(.A1(new_n733_), .A2(new_n797_), .ZN(new_n1307_));
  INV_X1    g0929(.A(new_n1086_), .ZN(new_n1308_));
  XNOR2_X1  g0930(.A(new_n1307_), .B(new_n1308_), .ZN(G324));
  XOR2_X1   g0931(.A(new_n1060_), .B(KEYINPUT39), .Z(G252));
  OAI21_X1  g0932(.A(new_n446_), .B1(new_n1091_), .B2(new_n494_), .ZN(G276));
  INV_X1    g0933(.A(KEYINPUT40), .ZN(new_n1312_));
  NAND2_X1  g0934(.A1(new_n563_), .A2(new_n1312_), .ZN(new_n1313_));
  NAND3_X1  g0935(.A1(new_n542_), .A2(KEYINPUT40), .A3(new_n562_), .ZN(new_n1314_));
  NAND2_X1  g0936(.A1(new_n1313_), .A2(new_n1314_), .ZN(new_n1315_));
  NAND2_X1  g0937(.A1(new_n1315_), .A2(new_n561_), .ZN(new_n1316_));
  INV_X1    g0938(.A(new_n1081_), .ZN(new_n1317_));
  INV_X1    g0939(.A(new_n586_), .ZN(new_n1318_));
  NOR2_X1   g0940(.A1(new_n1317_), .A2(new_n1318_), .ZN(new_n1319_));
  AOI21_X1  g0941(.A(G2224), .B1(new_n531_), .B2(new_n532_), .ZN(new_n1320_));
  OAI211_X1 g0942(.A(new_n532_), .B(G2224), .C1(G18), .C2(new_n529_), .ZN(new_n1321_));
  INV_X1    g0943(.A(new_n1321_), .ZN(new_n1322_));
  NOR2_X1   g0944(.A1(new_n1320_), .A2(new_n1322_), .ZN(new_n1323_));
  INV_X1    g0945(.A(new_n1323_), .ZN(new_n1324_));
  NOR2_X1   g0946(.A1(new_n1324_), .A2(new_n541_), .ZN(new_n1325_));
  AOI21_X1  g0947(.A(new_n1316_), .B1(new_n1319_), .B2(new_n1325_), .ZN(new_n1326_));
  XOR2_X1   g0948(.A(new_n1326_), .B(new_n588_), .Z(G310));
  INV_X1    g0949(.A(new_n562_), .ZN(new_n1328_));
  OAI21_X1  g0950(.A(new_n535_), .B1(new_n1328_), .B2(new_n1322_), .ZN(new_n1329_));
  AOI21_X1  g0951(.A(new_n1329_), .B1(new_n560_), .B2(new_n539_), .ZN(new_n1330_));
  INV_X1    g0952(.A(new_n1319_), .ZN(new_n1331_));
  OAI21_X1  g0953(.A(new_n1330_), .B1(new_n1331_), .B2(new_n540_), .ZN(new_n1332_));
  XNOR2_X1  g0954(.A(new_n1332_), .B(new_n541_), .ZN(G313));
  INV_X1    g0955(.A(new_n548_), .ZN(new_n1334_));
  OAI21_X1  g0956(.A(new_n558_), .B1(new_n1334_), .B2(new_n552_), .ZN(new_n1335_));
  NAND2_X1  g0957(.A1(new_n1335_), .A2(new_n1328_), .ZN(new_n1336_));
  NOR2_X1   g0958(.A1(new_n1319_), .A2(new_n1336_), .ZN(new_n1337_));
  XNOR2_X1  g0959(.A(new_n1337_), .B(new_n1323_), .ZN(G316));
  AOI21_X1  g0960(.A(new_n558_), .B1(new_n1081_), .B2(new_n584_), .ZN(new_n1339_));
  XOR2_X1   g0961(.A(new_n1339_), .B(new_n554_), .Z(G319));
  NOR2_X1   g0962(.A1(new_n482_), .A2(new_n470_), .ZN(new_n1341_));
  OAI21_X1  g0963(.A(new_n456_), .B1(new_n458_), .B2(new_n477_), .ZN(new_n1342_));
  AOI21_X1  g0964(.A(new_n1341_), .B1(new_n741_), .B2(new_n1342_), .ZN(new_n1343_));
  OAI21_X1  g0965(.A(new_n1308_), .B1(new_n733_), .B2(new_n797_), .ZN(new_n1344_));
  OAI21_X1  g0966(.A(new_n1343_), .B1(new_n1344_), .B2(new_n1085_), .ZN(new_n1345_));
  XNOR2_X1  g0967(.A(new_n1345_), .B(new_n466_), .ZN(G327));
  OAI21_X1  g0968(.A(KEYINPUT41), .B1(new_n483_), .B2(new_n456_), .ZN(new_n1347_));
  INV_X1    g0969(.A(KEYINPUT41), .ZN(new_n1348_));
  NAND4_X1  g0970(.A1(new_n457_), .A2(new_n449_), .A3(new_n1348_), .A4(new_n451_), .ZN(new_n1349_));
  AND3_X1   g0971(.A1(new_n1347_), .A2(new_n451_), .A3(new_n1349_), .ZN(new_n1350_));
  AND2_X1   g0972(.A1(new_n1344_), .A2(new_n477_), .ZN(new_n1351_));
  OAI21_X1  g0973(.A(new_n1350_), .B1(new_n1351_), .B2(new_n460_), .ZN(new_n1352_));
  XNOR2_X1  g0974(.A(new_n1352_), .B(new_n473_), .ZN(G330));
  INV_X1    g0975(.A(new_n1342_), .ZN(new_n1354_));
  OAI21_X1  g0976(.A(new_n1354_), .B1(new_n1307_), .B2(new_n740_), .ZN(new_n1355_));
  XNOR2_X1  g0977(.A(new_n1355_), .B(new_n483_), .ZN(G333));
  XNOR2_X1  g0978(.A(new_n1351_), .B(new_n459_), .ZN(G336));
  OR4_X1    g0979(.A1(G404), .A2(G406), .A3(G408), .A4(G410), .ZN(new_n1358_));
  NOR3_X1   g0980(.A1(G414), .A2(G416), .A3(new_n1358_), .ZN(new_n1359_));
  NAND3_X1  g0981(.A1(new_n1359_), .A2(new_n1198_), .A3(new_n1197_), .ZN(G418));
  INV_X1    g0982(.A(new_n740_), .ZN(new_n1361_));
  NOR2_X1   g0983(.A1(new_n742_), .A2(new_n466_), .ZN(new_n1362_));
  OAI211_X1 g0984(.A(new_n1361_), .B(new_n1362_), .C1(new_n733_), .C2(new_n797_), .ZN(new_n1363_));
  NAND2_X1  g0985(.A1(new_n1363_), .A2(new_n487_), .ZN(new_n1364_));
  INV_X1    g0986(.A(new_n1364_), .ZN(new_n1365_));
  OAI21_X1  g0987(.A(new_n446_), .B1(new_n1365_), .B2(new_n494_), .ZN(G273));
  AOI21_X1  g0988(.A(new_n571_), .B1(new_n1081_), .B2(new_n590_), .ZN(new_n1367_));
  INV_X1    g0989(.A(new_n521_), .ZN(new_n1368_));
  NAND2_X1  g0990(.A1(new_n1367_), .A2(new_n1368_), .ZN(new_n1369_));
  NAND2_X1  g0991(.A1(new_n509_), .A2(new_n576_), .ZN(new_n1370_));
  NAND2_X1  g0992(.A1(new_n1370_), .A2(new_n508_), .ZN(new_n1371_));
  AOI21_X1  g0993(.A(new_n504_), .B1(new_n1371_), .B2(new_n520_), .ZN(new_n1372_));
  OAI21_X1  g0994(.A(new_n1369_), .B1(new_n1367_), .B2(new_n1372_), .ZN(new_n1373_));
  XOR2_X1   g0995(.A(new_n1373_), .B(new_n579_), .Z(G298));
  NAND2_X1  g0996(.A1(new_n520_), .A2(new_n503_), .ZN(new_n1375_));
  XOR2_X1   g0997(.A(new_n1375_), .B(new_n517_), .Z(new_n1376_));
  AND3_X1   g0998(.A1(new_n1367_), .A2(KEYINPUT42), .A3(new_n1376_), .ZN(new_n1377_));
  AOI21_X1  g0999(.A(KEYINPUT42), .B1(new_n1367_), .B2(new_n1376_), .ZN(new_n1378_));
  XNOR2_X1  g1000(.A(new_n1375_), .B(new_n1371_), .ZN(new_n1379_));
  OR2_X1    g1001(.A1(new_n1367_), .A2(new_n1379_), .ZN(new_n1380_));
  AOI21_X1  g1002(.A(new_n1377_), .B1(new_n1378_), .B2(new_n1380_), .ZN(G301));
  OAI21_X1  g1003(.A(new_n515_), .B1(new_n1367_), .B2(new_n576_), .ZN(new_n1382_));
  INV_X1    g1004(.A(new_n574_), .ZN(new_n1383_));
  XNOR2_X1  g1005(.A(new_n1382_), .B(new_n1383_), .ZN(G304));
  XNOR2_X1  g1006(.A(new_n1367_), .B(new_n577_), .ZN(G307));
  INV_X1    g1007(.A(new_n1128_), .ZN(new_n1386_));
  NAND2_X1  g1008(.A1(new_n1386_), .A2(new_n619_), .ZN(new_n1387_));
  INV_X1    g1009(.A(new_n746_), .ZN(new_n1388_));
  NAND2_X1  g1010(.A1(new_n1387_), .A2(new_n1388_), .ZN(new_n1389_));
  INV_X1    g1011(.A(G4394), .ZN(new_n1390_));
  NAND2_X1  g1012(.A1(new_n1185_), .A2(new_n1390_), .ZN(new_n1391_));
  NAND2_X1  g1013(.A1(new_n1391_), .A2(new_n707_), .ZN(new_n1392_));
  XNOR2_X1  g1014(.A(new_n1389_), .B(new_n1392_), .ZN(G344));
  XNOR2_X1  g1015(.A(new_n493_), .B(new_n491_), .ZN(new_n1394_));
  NOR2_X1   g1016(.A1(new_n1364_), .A2(new_n1394_), .ZN(new_n1395_));
  INV_X1    g1017(.A(new_n1395_), .ZN(new_n1396_));
  AOI22_X1  g1018(.A1(new_n493_), .A2(new_n445_), .B1(new_n442_), .B2(new_n489_), .ZN(new_n1397_));
  OAI21_X1  g1019(.A(new_n1396_), .B1(new_n1365_), .B2(new_n1397_), .ZN(G422));
  INV_X1    g1020(.A(KEYINPUT43), .ZN(new_n1399_));
  OAI211_X1 g1021(.A(new_n1396_), .B(new_n1399_), .C1(new_n1365_), .C2(new_n1397_), .ZN(new_n1400_));
  NOR2_X1   g1022(.A1(new_n1365_), .A2(new_n1397_), .ZN(new_n1401_));
  OAI21_X1  g1023(.A(KEYINPUT43), .B1(new_n1401_), .B2(new_n1395_), .ZN(new_n1402_));
  NAND2_X1  g1024(.A1(new_n1400_), .A2(new_n1402_), .ZN(G469));
  XNOR2_X1  g1025(.A(new_n1364_), .B(new_n492_), .ZN(G419));
  XNOR2_X1  g1026(.A(new_n1364_), .B(new_n492_), .ZN(G471));
  NAND2_X1  g1027(.A1(new_n701_), .A2(new_n703_), .ZN(new_n1406_));
  NOR2_X1   g1028(.A1(new_n1406_), .A2(new_n1392_), .ZN(new_n1407_));
  NAND3_X1  g1029(.A1(new_n1389_), .A2(new_n1407_), .A3(new_n790_), .ZN(new_n1408_));
  NAND4_X1  g1030(.A1(new_n704_), .A2(new_n716_), .A3(new_n723_), .A4(new_n709_), .ZN(new_n1409_));
  AOI21_X1  g1031(.A(new_n720_), .B1(new_n701_), .B2(new_n788_), .ZN(new_n1410_));
  AOI21_X1  g1032(.A(new_n715_), .B1(new_n1410_), .B2(new_n713_), .ZN(new_n1411_));
  NAND3_X1  g1033(.A1(new_n1408_), .A2(new_n1409_), .A3(new_n1411_), .ZN(new_n1412_));
  XNOR2_X1  g1034(.A(new_n1412_), .B(new_n729_), .ZN(G359));
  AOI21_X1  g1035(.A(new_n792_), .B1(new_n1389_), .B2(new_n1407_), .ZN(new_n1414_));
  OAI21_X1  g1036(.A(new_n788_), .B1(new_n1414_), .B2(new_n720_), .ZN(new_n1415_));
  INV_X1    g1037(.A(new_n716_), .ZN(new_n1416_));
  XNOR2_X1  g1038(.A(new_n1415_), .B(new_n1416_), .ZN(G362));
  XNOR2_X1  g1039(.A(new_n1414_), .B(new_n723_), .ZN(G365));
  AOI21_X1  g1040(.A(new_n709_), .B1(new_n1389_), .B2(new_n707_), .ZN(new_n1419_));
  XNOR2_X1  g1041(.A(new_n1419_), .B(new_n704_), .ZN(G368));
  INV_X1    g1042(.A(new_n794_), .ZN(new_n1421_));
  OAI21_X1  g1043(.A(new_n1421_), .B1(new_n1408_), .B2(new_n729_), .ZN(new_n1422_));
  NAND3_X1  g1044(.A1(new_n772_), .A2(new_n695_), .A3(new_n688_), .ZN(new_n1423_));
  NAND2_X1  g1045(.A1(new_n775_), .A2(new_n1423_), .ZN(new_n1424_));
  XNOR2_X1  g1046(.A(new_n1424_), .B(KEYINPUT44), .ZN(new_n1425_));
  NOR2_X1   g1047(.A1(new_n1422_), .A2(new_n1425_), .ZN(new_n1426_));
  NOR2_X1   g1048(.A1(new_n672_), .A2(new_n680_), .ZN(new_n1427_));
  INV_X1    g1049(.A(new_n1427_), .ZN(new_n1428_));
  OAI211_X1 g1050(.A(new_n689_), .B(new_n1428_), .C1(new_n675_), .C2(new_n672_), .ZN(new_n1429_));
  NAND2_X1  g1051(.A1(new_n1429_), .A2(new_n688_), .ZN(new_n1430_));
  XNOR2_X1  g1052(.A(new_n1430_), .B(new_n774_), .ZN(new_n1431_));
  AOI21_X1  g1053(.A(new_n1426_), .B1(new_n1422_), .B2(new_n1431_), .ZN(G347));
  AOI21_X1  g1054(.A(new_n682_), .B1(new_n1422_), .B2(new_n680_), .ZN(new_n1433_));
  INV_X1    g1055(.A(new_n675_), .ZN(new_n1434_));
  OAI21_X1  g1056(.A(new_n664_), .B1(new_n1433_), .B2(new_n1434_), .ZN(new_n1435_));
  XNOR2_X1  g1057(.A(new_n1435_), .B(new_n690_), .ZN(G350));
  XNOR2_X1  g1058(.A(new_n1433_), .B(new_n675_), .ZN(G353));
  INV_X1    g1059(.A(new_n683_), .ZN(new_n1438_));
  XNOR2_X1  g1060(.A(new_n1422_), .B(new_n1438_), .ZN(G356));
  AOI21_X1  g1061(.A(new_n1316_), .B1(new_n542_), .B2(new_n586_), .ZN(new_n1440_));
  NAND2_X1  g1062(.A1(new_n1305_), .A2(new_n554_), .ZN(new_n1441_));
  OAI21_X1  g1063(.A(KEYINPUT47), .B1(new_n586_), .B2(new_n1336_), .ZN(new_n1442_));
  INV_X1    g1064(.A(new_n1442_), .ZN(new_n1443_));
  NOR3_X1   g1065(.A1(new_n586_), .A2(new_n1336_), .A3(KEYINPUT47), .ZN(new_n1444_));
  OAI211_X1 g1066(.A(new_n1318_), .B(new_n1441_), .C1(new_n1443_), .C2(new_n1444_), .ZN(new_n1445_));
  NOR2_X1   g1067(.A1(new_n554_), .A2(new_n585_), .ZN(new_n1446_));
  AOI21_X1  g1068(.A(new_n1329_), .B1(new_n1446_), .B2(new_n539_), .ZN(new_n1447_));
  INV_X1    g1069(.A(new_n1444_), .ZN(new_n1448_));
  NAND2_X1  g1070(.A1(new_n1318_), .A2(new_n1441_), .ZN(new_n1449_));
  NAND3_X1  g1071(.A1(new_n1448_), .A2(new_n1449_), .A3(new_n1442_), .ZN(new_n1450_));
  AND3_X1   g1072(.A1(new_n1445_), .A2(new_n1447_), .A3(new_n1450_), .ZN(new_n1451_));
  AOI21_X1  g1073(.A(new_n1447_), .B1(new_n1445_), .B2(new_n1450_), .ZN(new_n1452_));
  OAI21_X1  g1074(.A(new_n1440_), .B1(new_n1451_), .B2(new_n1452_), .ZN(new_n1453_));
  NAND2_X1  g1075(.A1(new_n1445_), .A2(new_n1450_), .ZN(new_n1454_));
  INV_X1    g1076(.A(new_n1447_), .ZN(new_n1455_));
  NAND2_X1  g1077(.A1(new_n1454_), .A2(new_n1455_), .ZN(new_n1456_));
  INV_X1    g1078(.A(new_n1316_), .ZN(new_n1457_));
  NAND2_X1  g1079(.A1(new_n1457_), .A2(new_n587_), .ZN(new_n1458_));
  NAND3_X1  g1080(.A1(new_n1445_), .A2(new_n1447_), .A3(new_n1450_), .ZN(new_n1459_));
  NAND3_X1  g1081(.A1(new_n1456_), .A2(new_n1458_), .A3(new_n1459_), .ZN(new_n1460_));
  OR2_X1    g1082(.A1(new_n585_), .A2(KEYINPUT46), .ZN(new_n1461_));
  XNOR2_X1  g1083(.A(new_n588_), .B(new_n1461_), .ZN(new_n1462_));
  AND3_X1   g1084(.A1(new_n1453_), .A2(new_n1460_), .A3(new_n1462_), .ZN(new_n1463_));
  AOI21_X1  g1085(.A(new_n1462_), .B1(new_n1453_), .B2(new_n1460_), .ZN(new_n1464_));
  OAI21_X1  g1086(.A(new_n1323_), .B1(new_n1463_), .B2(new_n1464_), .ZN(new_n1465_));
  INV_X1    g1087(.A(new_n1462_), .ZN(new_n1466_));
  NOR3_X1   g1088(.A1(new_n1451_), .A2(new_n1440_), .A3(new_n1452_), .ZN(new_n1467_));
  AOI21_X1  g1089(.A(new_n1458_), .B1(new_n1456_), .B2(new_n1459_), .ZN(new_n1468_));
  OAI21_X1  g1090(.A(new_n1466_), .B1(new_n1467_), .B2(new_n1468_), .ZN(new_n1469_));
  NAND3_X1  g1091(.A1(new_n1453_), .A2(new_n1460_), .A3(new_n1462_), .ZN(new_n1470_));
  NAND3_X1  g1092(.A1(new_n1469_), .A2(new_n540_), .A3(new_n1470_), .ZN(new_n1471_));
  AND3_X1   g1093(.A1(new_n1465_), .A2(new_n541_), .A3(new_n1471_), .ZN(new_n1472_));
  AOI21_X1  g1094(.A(new_n541_), .B1(new_n1465_), .B2(new_n1471_), .ZN(new_n1473_));
  OAI21_X1  g1095(.A(new_n1081_), .B1(new_n1472_), .B2(new_n1473_), .ZN(new_n1474_));
  NAND2_X1  g1096(.A1(new_n1329_), .A2(new_n559_), .ZN(new_n1475_));
  OAI211_X1 g1097(.A(new_n535_), .B(new_n558_), .C1(new_n1328_), .C2(new_n1322_), .ZN(new_n1476_));
  INV_X1    g1098(.A(new_n1335_), .ZN(new_n1477_));
  AOI22_X1  g1099(.A1(new_n1475_), .A2(new_n1476_), .B1(new_n1477_), .B2(new_n1321_), .ZN(new_n1478_));
  OR2_X1    g1100(.A1(new_n1449_), .A2(new_n1478_), .ZN(new_n1479_));
  NAND2_X1  g1101(.A1(new_n1449_), .A2(new_n1478_), .ZN(new_n1480_));
  NAND2_X1  g1102(.A1(new_n1479_), .A2(new_n1480_), .ZN(new_n1481_));
  NAND2_X1  g1103(.A1(new_n1457_), .A2(new_n1481_), .ZN(new_n1482_));
  XNOR2_X1  g1104(.A(new_n588_), .B(new_n1336_), .ZN(new_n1483_));
  NAND3_X1  g1105(.A1(new_n1316_), .A2(new_n1479_), .A3(new_n1480_), .ZN(new_n1484_));
  NAND3_X1  g1106(.A1(new_n1482_), .A2(new_n1483_), .A3(new_n1484_), .ZN(new_n1485_));
  INV_X1    g1107(.A(new_n1485_), .ZN(new_n1486_));
  AOI21_X1  g1108(.A(new_n1483_), .B1(new_n1482_), .B2(new_n1484_), .ZN(new_n1487_));
  OAI21_X1  g1109(.A(new_n540_), .B1(new_n1486_), .B2(new_n1487_), .ZN(new_n1488_));
  OR2_X1    g1110(.A1(new_n541_), .A2(KEYINPUT48), .ZN(new_n1489_));
  NAND2_X1  g1111(.A1(new_n1482_), .A2(new_n1484_), .ZN(new_n1490_));
  INV_X1    g1112(.A(new_n1483_), .ZN(new_n1491_));
  NAND2_X1  g1113(.A1(new_n1490_), .A2(new_n1491_), .ZN(new_n1492_));
  NAND3_X1  g1114(.A1(new_n1492_), .A2(new_n1323_), .A3(new_n1485_), .ZN(new_n1493_));
  NAND3_X1  g1115(.A1(new_n1488_), .A2(new_n1489_), .A3(new_n1493_), .ZN(new_n1494_));
  NAND3_X1  g1116(.A1(new_n1494_), .A2(KEYINPUT48), .A3(new_n541_), .ZN(new_n1495_));
  NAND2_X1  g1117(.A1(new_n541_), .A2(KEYINPUT48), .ZN(new_n1496_));
  NAND4_X1  g1118(.A1(new_n1488_), .A2(new_n1493_), .A3(new_n1496_), .A4(new_n1489_), .ZN(new_n1497_));
  NAND2_X1  g1119(.A1(new_n1495_), .A2(new_n1497_), .ZN(new_n1498_));
  OR2_X1    g1120(.A1(new_n1081_), .A2(KEYINPUT45), .ZN(new_n1499_));
  NAND2_X1  g1121(.A1(new_n1081_), .A2(KEYINPUT45), .ZN(new_n1500_));
  NAND2_X1  g1122(.A1(new_n1499_), .A2(new_n1500_), .ZN(new_n1501_));
  INV_X1    g1123(.A(new_n1501_), .ZN(new_n1502_));
  NAND2_X1  g1124(.A1(new_n1498_), .A2(new_n1502_), .ZN(new_n1503_));
  NAND2_X1  g1125(.A1(new_n1474_), .A2(new_n1503_), .ZN(new_n1504_));
  INV_X1    g1126(.A(new_n1370_), .ZN(new_n1505_));
  NOR2_X1   g1127(.A1(new_n509_), .A2(new_n576_), .ZN(new_n1506_));
  OAI21_X1  g1128(.A(new_n515_), .B1(new_n1505_), .B2(new_n1506_), .ZN(new_n1507_));
  OAI21_X1  g1129(.A(new_n1507_), .B1(new_n573_), .B2(new_n515_), .ZN(new_n1508_));
  XNOR2_X1  g1130(.A(new_n1508_), .B(new_n579_), .ZN(new_n1509_));
  OR2_X1    g1131(.A1(new_n1509_), .A2(new_n1368_), .ZN(new_n1510_));
  NAND2_X1  g1132(.A1(new_n1509_), .A2(new_n1368_), .ZN(new_n1511_));
  NAND2_X1  g1133(.A1(new_n1510_), .A2(new_n1511_), .ZN(new_n1512_));
  NAND2_X1  g1134(.A1(new_n1383_), .A2(new_n1375_), .ZN(new_n1513_));
  AND2_X1   g1135(.A1(new_n1513_), .A2(new_n575_), .ZN(new_n1514_));
  INV_X1    g1136(.A(new_n1514_), .ZN(new_n1515_));
  XNOR2_X1  g1137(.A(new_n1512_), .B(new_n1515_), .ZN(new_n1516_));
  NAND2_X1  g1138(.A1(new_n1516_), .A2(new_n572_), .ZN(new_n1517_));
  XNOR2_X1  g1139(.A(new_n508_), .B(new_n515_), .ZN(new_n1518_));
  OAI21_X1  g1140(.A(new_n1370_), .B1(new_n1518_), .B2(new_n576_), .ZN(new_n1519_));
  XOR2_X1   g1141(.A(new_n1519_), .B(new_n579_), .Z(new_n1520_));
  NAND2_X1  g1142(.A1(new_n1520_), .A2(new_n574_), .ZN(new_n1521_));
  XNOR2_X1  g1143(.A(new_n1519_), .B(new_n579_), .ZN(new_n1522_));
  NAND2_X1  g1144(.A1(new_n1522_), .A2(new_n1383_), .ZN(new_n1523_));
  NAND2_X1  g1145(.A1(new_n1521_), .A2(new_n1523_), .ZN(new_n1524_));
  INV_X1    g1146(.A(new_n520_), .ZN(new_n1525_));
  AOI21_X1  g1147(.A(new_n1525_), .B1(new_n503_), .B2(new_n1371_), .ZN(new_n1526_));
  INV_X1    g1148(.A(new_n1526_), .ZN(new_n1527_));
  NAND2_X1  g1149(.A1(new_n1524_), .A2(new_n1527_), .ZN(new_n1528_));
  NAND3_X1  g1150(.A1(new_n1521_), .A2(new_n1526_), .A3(new_n1523_), .ZN(new_n1529_));
  AND2_X1   g1151(.A1(new_n1528_), .A2(new_n1529_), .ZN(new_n1530_));
  OAI211_X1 g1152(.A(new_n1502_), .B(new_n1517_), .C1(new_n572_), .C2(new_n1530_), .ZN(new_n1531_));
  AND2_X1   g1153(.A1(new_n572_), .A2(new_n589_), .ZN(new_n1532_));
  NAND2_X1  g1154(.A1(new_n1516_), .A2(new_n1532_), .ZN(new_n1533_));
  OAI211_X1 g1155(.A(new_n1533_), .B(new_n1081_), .C1(new_n1532_), .C2(new_n1530_), .ZN(new_n1534_));
  AND2_X1   g1156(.A1(new_n1531_), .A2(new_n1534_), .ZN(new_n1535_));
  NAND3_X1  g1157(.A1(new_n1469_), .A2(new_n1324_), .A3(new_n1470_), .ZN(new_n1536_));
  NAND2_X1  g1158(.A1(new_n1536_), .A2(new_n541_), .ZN(new_n1537_));
  AOI21_X1  g1159(.A(new_n540_), .B1(new_n1469_), .B2(new_n1470_), .ZN(new_n1538_));
  NOR2_X1   g1160(.A1(new_n1537_), .A2(new_n1538_), .ZN(new_n1539_));
  OAI21_X1  g1161(.A(new_n1501_), .B1(new_n1539_), .B2(new_n1473_), .ZN(new_n1540_));
  AOI22_X1  g1162(.A1(new_n1498_), .A2(new_n1317_), .B1(new_n1531_), .B2(new_n1534_), .ZN(new_n1541_));
  AOI22_X1  g1163(.A1(new_n1504_), .A2(new_n1535_), .B1(new_n1540_), .B2(new_n1541_), .ZN(G321));
  OAI21_X1  g1164(.A(new_n1342_), .B1(new_n741_), .B2(new_n1341_), .ZN(new_n1543_));
  OAI21_X1  g1165(.A(new_n1543_), .B1(new_n1342_), .B2(new_n1341_), .ZN(new_n1544_));
  INV_X1    g1166(.A(new_n1544_), .ZN(new_n1545_));
  NAND2_X1  g1167(.A1(new_n1350_), .A2(new_n477_), .ZN(new_n1546_));
  NAND4_X1  g1168(.A1(new_n460_), .A2(new_n1347_), .A3(new_n451_), .A4(new_n1349_), .ZN(new_n1547_));
  INV_X1    g1169(.A(new_n477_), .ZN(new_n1548_));
  NAND2_X1  g1170(.A1(new_n1547_), .A2(new_n1548_), .ZN(new_n1549_));
  NAND3_X1  g1171(.A1(new_n1546_), .A2(new_n1549_), .A3(new_n1086_), .ZN(new_n1550_));
  INV_X1    g1172(.A(new_n1550_), .ZN(new_n1551_));
  AOI21_X1  g1173(.A(new_n1086_), .B1(new_n1546_), .B2(new_n1549_), .ZN(new_n1552_));
  OAI21_X1  g1174(.A(new_n1545_), .B1(new_n1551_), .B2(new_n1552_), .ZN(new_n1553_));
  NAND2_X1  g1175(.A1(new_n1546_), .A2(new_n1549_), .ZN(new_n1554_));
  NAND2_X1  g1176(.A1(new_n1554_), .A2(new_n1308_), .ZN(new_n1555_));
  NAND3_X1  g1177(.A1(new_n1555_), .A2(new_n1550_), .A3(new_n1544_), .ZN(new_n1556_));
  NAND3_X1  g1178(.A1(new_n1553_), .A2(new_n1556_), .A3(new_n1084_), .ZN(new_n1557_));
  AOI21_X1  g1179(.A(new_n459_), .B1(new_n1553_), .B2(new_n1556_), .ZN(new_n1558_));
  OAI21_X1  g1180(.A(new_n1557_), .B1(new_n1558_), .B2(KEYINPUT51), .ZN(new_n1559_));
  INV_X1    g1181(.A(KEYINPUT51), .ZN(new_n1560_));
  AOI211_X1 g1182(.A(new_n1560_), .B(new_n459_), .C1(new_n1553_), .C2(new_n1556_), .ZN(new_n1561_));
  OAI21_X1  g1183(.A(new_n466_), .B1(new_n1559_), .B2(new_n1561_), .ZN(new_n1562_));
  NOR3_X1   g1184(.A1(new_n1551_), .A2(new_n1552_), .A3(new_n1545_), .ZN(new_n1563_));
  AOI21_X1  g1185(.A(new_n1544_), .B1(new_n1555_), .B2(new_n1550_), .ZN(new_n1564_));
  OAI21_X1  g1186(.A(new_n1084_), .B1(new_n1563_), .B2(new_n1564_), .ZN(new_n1565_));
  INV_X1    g1187(.A(new_n459_), .ZN(new_n1566_));
  NAND3_X1  g1188(.A1(new_n1553_), .A2(new_n1556_), .A3(new_n1566_), .ZN(new_n1567_));
  AOI21_X1  g1189(.A(new_n466_), .B1(new_n1565_), .B2(new_n1567_), .ZN(new_n1568_));
  INV_X1    g1190(.A(new_n1568_), .ZN(new_n1569_));
  AOI21_X1  g1191(.A(new_n483_), .B1(new_n1562_), .B2(new_n1569_), .ZN(new_n1570_));
  NAND3_X1  g1192(.A1(new_n1565_), .A2(new_n466_), .A3(new_n1567_), .ZN(new_n1571_));
  AND3_X1   g1193(.A1(new_n1569_), .A2(new_n1571_), .A3(new_n483_), .ZN(new_n1572_));
  OAI21_X1  g1194(.A(new_n473_), .B1(new_n1570_), .B2(new_n1572_), .ZN(new_n1573_));
  INV_X1    g1195(.A(new_n473_), .ZN(new_n1574_));
  NAND3_X1  g1196(.A1(new_n1569_), .A2(new_n1571_), .A3(new_n483_), .ZN(new_n1575_));
  OAI21_X1  g1197(.A(new_n1566_), .B1(new_n1563_), .B2(new_n1564_), .ZN(new_n1576_));
  NAND2_X1  g1198(.A1(new_n1576_), .A2(new_n1560_), .ZN(new_n1577_));
  NAND2_X1  g1199(.A1(new_n1558_), .A2(KEYINPUT51), .ZN(new_n1578_));
  NAND3_X1  g1200(.A1(new_n1577_), .A2(new_n1578_), .A3(new_n1557_), .ZN(new_n1579_));
  AOI21_X1  g1201(.A(new_n1568_), .B1(new_n1579_), .B2(new_n466_), .ZN(new_n1580_));
  OAI211_X1 g1202(.A(new_n1574_), .B(new_n1575_), .C1(new_n1580_), .C2(new_n483_), .ZN(new_n1581_));
  NAND2_X1  g1203(.A1(new_n1573_), .A2(new_n1581_), .ZN(new_n1582_));
  NAND2_X1  g1204(.A1(new_n1582_), .A2(new_n1083_), .ZN(new_n1583_));
  INV_X1    g1205(.A(new_n466_), .ZN(new_n1584_));
  NAND2_X1  g1206(.A1(new_n740_), .A2(new_n1354_), .ZN(new_n1585_));
  NAND2_X1  g1207(.A1(new_n1585_), .A2(new_n1341_), .ZN(new_n1586_));
  AOI21_X1  g1208(.A(new_n741_), .B1(new_n740_), .B2(new_n1354_), .ZN(new_n1587_));
  OR2_X1    g1209(.A1(new_n1587_), .A2(new_n1341_), .ZN(new_n1588_));
  NAND2_X1  g1210(.A1(new_n1547_), .A2(new_n737_), .ZN(new_n1589_));
  NOR2_X1   g1211(.A1(new_n1589_), .A2(new_n1308_), .ZN(new_n1590_));
  NAND4_X1  g1212(.A1(new_n1347_), .A2(new_n739_), .A3(new_n451_), .A4(new_n1349_), .ZN(new_n1591_));
  AOI21_X1  g1213(.A(new_n1591_), .B1(new_n1547_), .B2(new_n737_), .ZN(new_n1592_));
  OAI211_X1 g1214(.A(new_n1586_), .B(new_n1588_), .C1(new_n1590_), .C2(new_n1592_), .ZN(new_n1593_));
  OAI21_X1  g1215(.A(new_n1586_), .B1(new_n1341_), .B2(new_n1587_), .ZN(new_n1594_));
  INV_X1    g1216(.A(new_n737_), .ZN(new_n1595_));
  OAI211_X1 g1217(.A(new_n1350_), .B(new_n739_), .C1(new_n1595_), .C2(new_n460_), .ZN(new_n1596_));
  OAI211_X1 g1218(.A(new_n1594_), .B(new_n1596_), .C1(new_n1308_), .C2(new_n1589_), .ZN(new_n1597_));
  AND3_X1   g1219(.A1(new_n1593_), .A2(new_n1597_), .A3(new_n1084_), .ZN(new_n1598_));
  AOI21_X1  g1220(.A(new_n459_), .B1(new_n1593_), .B2(new_n1597_), .ZN(new_n1599_));
  OAI21_X1  g1221(.A(new_n1584_), .B1(new_n1598_), .B2(new_n1599_), .ZN(new_n1600_));
  NAND2_X1  g1222(.A1(new_n1593_), .A2(new_n1597_), .ZN(new_n1601_));
  NAND2_X1  g1223(.A1(new_n1601_), .A2(new_n1566_), .ZN(new_n1602_));
  NAND3_X1  g1224(.A1(new_n1593_), .A2(new_n1597_), .A3(new_n1084_), .ZN(new_n1603_));
  NAND3_X1  g1225(.A1(new_n1602_), .A2(new_n466_), .A3(new_n1603_), .ZN(new_n1604_));
  NAND3_X1  g1226(.A1(new_n1600_), .A2(new_n1604_), .A3(KEYINPUT49), .ZN(new_n1605_));
  INV_X1    g1227(.A(KEYINPUT49), .ZN(new_n1606_));
  NAND4_X1  g1228(.A1(new_n1602_), .A2(new_n1606_), .A3(new_n466_), .A4(new_n1603_), .ZN(new_n1607_));
  NAND3_X1  g1229(.A1(new_n1605_), .A2(new_n483_), .A3(new_n1607_), .ZN(new_n1608_));
  INV_X1    g1230(.A(new_n1084_), .ZN(new_n1609_));
  AOI21_X1  g1231(.A(new_n1584_), .B1(new_n1601_), .B2(new_n1609_), .ZN(new_n1610_));
  OAI21_X1  g1232(.A(new_n1610_), .B1(new_n1566_), .B2(new_n1601_), .ZN(new_n1611_));
  NAND3_X1  g1233(.A1(new_n1611_), .A2(new_n452_), .A3(new_n1600_), .ZN(new_n1612_));
  NAND2_X1  g1234(.A1(new_n1608_), .A2(new_n1612_), .ZN(new_n1613_));
  NOR2_X1   g1235(.A1(new_n1613_), .A2(new_n473_), .ZN(new_n1614_));
  INV_X1    g1236(.A(KEYINPUT53), .ZN(new_n1615_));
  AOI21_X1  g1237(.A(new_n1574_), .B1(new_n1608_), .B2(new_n1612_), .ZN(new_n1616_));
  NOR3_X1   g1238(.A1(new_n1614_), .A2(new_n1615_), .A3(new_n1616_), .ZN(new_n1617_));
  INV_X1    g1239(.A(new_n1083_), .ZN(new_n1618_));
  INV_X1    g1240(.A(new_n1616_), .ZN(new_n1619_));
  OAI21_X1  g1241(.A(new_n1618_), .B1(new_n1619_), .B2(KEYINPUT53), .ZN(new_n1620_));
  OAI21_X1  g1242(.A(new_n1583_), .B1(new_n1617_), .B2(new_n1620_), .ZN(new_n1621_));
  XOR2_X1   g1243(.A(new_n1394_), .B(KEYINPUT52), .Z(new_n1622_));
  NAND2_X1  g1244(.A1(new_n1090_), .A2(new_n1622_), .ZN(new_n1623_));
  INV_X1    g1245(.A(new_n1397_), .ZN(new_n1624_));
  OAI211_X1 g1246(.A(new_n487_), .B(new_n1624_), .C1(new_n1083_), .C2(new_n1089_), .ZN(new_n1625_));
  AND2_X1   g1247(.A1(new_n1623_), .A2(new_n1625_), .ZN(new_n1626_));
  AOI21_X1  g1248(.A(new_n452_), .B1(new_n1611_), .B2(new_n1600_), .ZN(new_n1627_));
  NAND2_X1  g1249(.A1(new_n1605_), .A2(new_n1607_), .ZN(new_n1628_));
  NAND2_X1  g1250(.A1(new_n1628_), .A2(new_n452_), .ZN(new_n1629_));
  AOI21_X1  g1251(.A(new_n1627_), .B1(new_n1629_), .B2(KEYINPUT50), .ZN(new_n1630_));
  INV_X1    g1252(.A(KEYINPUT50), .ZN(new_n1631_));
  NAND3_X1  g1253(.A1(new_n1628_), .A2(new_n1631_), .A3(new_n452_), .ZN(new_n1632_));
  AOI21_X1  g1254(.A(new_n1574_), .B1(new_n1630_), .B2(new_n1632_), .ZN(new_n1633_));
  OAI21_X1  g1255(.A(new_n1618_), .B1(new_n1633_), .B2(new_n1614_), .ZN(new_n1634_));
  AOI21_X1  g1256(.A(new_n1626_), .B1(new_n1083_), .B2(new_n1582_), .ZN(new_n1635_));
  AOI22_X1  g1257(.A1(new_n1621_), .A2(new_n1626_), .B1(new_n1634_), .B2(new_n1635_), .ZN(G338));
  AOI21_X1  g1258(.A(G4400), .B1(new_n702_), .B2(new_n697_), .ZN(new_n1637_));
  OAI211_X1 g1259(.A(new_n713_), .B(new_n719_), .C1(new_n1637_), .C2(new_n722_), .ZN(new_n1638_));
  OAI211_X1 g1260(.A(new_n1638_), .B(new_n780_), .C1(new_n789_), .C2(new_n791_), .ZN(new_n1639_));
  MUX2_X1   g1261(.A(new_n1411_), .B(new_n1639_), .S(new_n792_), .Z(new_n1640_));
  XNOR2_X1  g1262(.A(new_n1640_), .B(new_n704_), .ZN(new_n1641_));
  XNOR2_X1  g1263(.A(new_n1641_), .B(new_n729_), .ZN(new_n1642_));
  INV_X1    g1264(.A(new_n723_), .ZN(new_n1643_));
  NAND2_X1  g1265(.A1(new_n1416_), .A2(new_n1643_), .ZN(new_n1644_));
  NAND2_X1  g1266(.A1(new_n1644_), .A2(new_n789_), .ZN(new_n1645_));
  XNOR2_X1  g1267(.A(new_n1642_), .B(new_n1645_), .ZN(new_n1646_));
  OAI21_X1  g1268(.A(new_n719_), .B1(new_n1637_), .B2(new_n722_), .ZN(new_n1647_));
  NAND3_X1  g1269(.A1(new_n701_), .A2(new_n703_), .A3(new_n719_), .ZN(new_n1648_));
  AOI21_X1  g1270(.A(new_n1391_), .B1(new_n1647_), .B2(new_n1648_), .ZN(new_n1649_));
  NOR2_X1   g1271(.A1(new_n1410_), .A2(new_n708_), .ZN(new_n1650_));
  INV_X1    g1272(.A(new_n1650_), .ZN(new_n1651_));
  NAND2_X1  g1273(.A1(new_n1410_), .A2(new_n708_), .ZN(new_n1652_));
  AOI21_X1  g1274(.A(new_n1649_), .B1(new_n1651_), .B2(new_n1652_), .ZN(new_n1653_));
  OR2_X1    g1275(.A1(new_n1646_), .A2(new_n1653_), .ZN(new_n1654_));
  INV_X1    g1276(.A(new_n1389_), .ZN(new_n1655_));
  NAND2_X1  g1277(.A1(new_n1646_), .A2(new_n1653_), .ZN(new_n1656_));
  NAND3_X1  g1278(.A1(new_n1654_), .A2(new_n1655_), .A3(new_n1656_), .ZN(new_n1657_));
  NOR2_X1   g1279(.A1(new_n1407_), .A2(new_n792_), .ZN(new_n1658_));
  XNOR2_X1  g1280(.A(new_n1658_), .B(new_n1392_), .ZN(new_n1659_));
  NAND2_X1  g1281(.A1(new_n788_), .A2(new_n707_), .ZN(new_n1660_));
  OAI21_X1  g1282(.A(new_n1647_), .B1(new_n1648_), .B2(new_n1660_), .ZN(new_n1661_));
  INV_X1    g1283(.A(new_n1661_), .ZN(new_n1662_));
  NOR3_X1   g1284(.A1(new_n789_), .A2(new_n1406_), .A3(new_n1392_), .ZN(new_n1663_));
  OAI21_X1  g1285(.A(new_n1662_), .B1(new_n1639_), .B2(new_n1663_), .ZN(new_n1664_));
  NAND4_X1  g1286(.A1(new_n1411_), .A2(new_n724_), .A3(new_n1409_), .A4(new_n1661_), .ZN(new_n1665_));
  NOR2_X1   g1287(.A1(new_n708_), .A2(KEYINPUT54), .ZN(new_n1666_));
  INV_X1    g1288(.A(new_n1666_), .ZN(new_n1667_));
  AND3_X1   g1289(.A1(new_n1664_), .A2(new_n1665_), .A3(new_n1667_), .ZN(new_n1668_));
  AOI21_X1  g1290(.A(new_n1667_), .B1(new_n1664_), .B2(new_n1665_), .ZN(new_n1669_));
  OAI21_X1  g1291(.A(new_n1659_), .B1(new_n1668_), .B2(new_n1669_), .ZN(new_n1670_));
  NAND2_X1  g1292(.A1(new_n1664_), .A2(new_n1665_), .ZN(new_n1671_));
  NAND2_X1  g1293(.A1(new_n1671_), .A2(new_n1666_), .ZN(new_n1672_));
  XNOR2_X1  g1294(.A(new_n1658_), .B(new_n710_), .ZN(new_n1673_));
  NAND3_X1  g1295(.A1(new_n1664_), .A2(new_n1665_), .A3(new_n1667_), .ZN(new_n1674_));
  NAND3_X1  g1296(.A1(new_n1672_), .A2(new_n1673_), .A3(new_n1674_), .ZN(new_n1675_));
  AND3_X1   g1297(.A1(new_n1670_), .A2(new_n1675_), .A3(new_n704_), .ZN(new_n1676_));
  AOI21_X1  g1298(.A(new_n704_), .B1(new_n1670_), .B2(new_n1675_), .ZN(new_n1677_));
  OAI21_X1  g1299(.A(new_n785_), .B1(new_n1676_), .B2(new_n1677_), .ZN(new_n1678_));
  NOR3_X1   g1300(.A1(new_n1668_), .A2(new_n1669_), .A3(new_n1659_), .ZN(new_n1679_));
  AOI21_X1  g1301(.A(new_n1673_), .B1(new_n1672_), .B2(new_n1674_), .ZN(new_n1680_));
  OAI21_X1  g1302(.A(new_n1406_), .B1(new_n1679_), .B2(new_n1680_), .ZN(new_n1681_));
  NAND3_X1  g1303(.A1(new_n1670_), .A2(new_n1675_), .A3(new_n704_), .ZN(new_n1682_));
  NAND3_X1  g1304(.A1(new_n1681_), .A2(new_n729_), .A3(new_n1682_), .ZN(new_n1683_));
  INV_X1    g1305(.A(KEYINPUT55), .ZN(new_n1684_));
  NAND3_X1  g1306(.A1(new_n1681_), .A2(new_n1684_), .A3(new_n729_), .ZN(new_n1685_));
  NAND3_X1  g1307(.A1(new_n1678_), .A2(new_n1683_), .A3(new_n1685_), .ZN(new_n1686_));
  NAND4_X1  g1308(.A1(new_n1681_), .A2(new_n1684_), .A3(new_n729_), .A4(new_n1682_), .ZN(new_n1687_));
  NAND3_X1  g1309(.A1(new_n1686_), .A2(new_n723_), .A3(new_n1687_), .ZN(new_n1688_));
  INV_X1    g1310(.A(KEYINPUT56), .ZN(new_n1689_));
  NAND4_X1  g1311(.A1(new_n1678_), .A2(new_n1683_), .A3(new_n1689_), .A4(new_n1643_), .ZN(new_n1690_));
  NAND3_X1  g1312(.A1(new_n1678_), .A2(new_n1683_), .A3(new_n1643_), .ZN(new_n1691_));
  NAND2_X1  g1313(.A1(new_n1691_), .A2(KEYINPUT56), .ZN(new_n1692_));
  NAND3_X1  g1314(.A1(new_n1688_), .A2(new_n1690_), .A3(new_n1692_), .ZN(new_n1693_));
  XNOR2_X1  g1315(.A(new_n1693_), .B(new_n716_), .ZN(new_n1694_));
  OAI21_X1  g1316(.A(new_n1657_), .B1(new_n1694_), .B2(new_n1655_), .ZN(new_n1695_));
  XNOR2_X1  g1317(.A(new_n675_), .B(new_n1438_), .ZN(new_n1696_));
  INV_X1    g1318(.A(new_n1696_), .ZN(new_n1697_));
  INV_X1    g1319(.A(new_n690_), .ZN(new_n1698_));
  INV_X1    g1320(.A(new_n1423_), .ZN(new_n1699_));
  AOI21_X1  g1321(.A(new_n695_), .B1(new_n772_), .B2(new_n688_), .ZN(new_n1700_));
  OAI21_X1  g1322(.A(new_n1698_), .B1(new_n1699_), .B2(new_n1700_), .ZN(new_n1701_));
  NAND3_X1  g1323(.A1(new_n775_), .A2(new_n690_), .A3(new_n1423_), .ZN(new_n1702_));
  NAND2_X1  g1324(.A1(new_n682_), .A2(new_n665_), .ZN(new_n1703_));
  NAND2_X1  g1325(.A1(new_n771_), .A2(new_n1703_), .ZN(new_n1704_));
  INV_X1    g1326(.A(new_n1704_), .ZN(new_n1705_));
  AND3_X1   g1327(.A1(new_n1701_), .A2(new_n1702_), .A3(new_n1705_), .ZN(new_n1706_));
  AOI21_X1  g1328(.A(new_n1705_), .B1(new_n1701_), .B2(new_n1702_), .ZN(new_n1707_));
  OAI21_X1  g1329(.A(new_n1697_), .B1(new_n1706_), .B2(new_n1707_), .ZN(new_n1708_));
  NAND2_X1  g1330(.A1(new_n1701_), .A2(new_n1702_), .ZN(new_n1709_));
  NAND2_X1  g1331(.A1(new_n1709_), .A2(new_n1704_), .ZN(new_n1710_));
  NAND3_X1  g1332(.A1(new_n1701_), .A2(new_n1702_), .A3(new_n1705_), .ZN(new_n1711_));
  NAND3_X1  g1333(.A1(new_n1710_), .A2(new_n1696_), .A3(new_n1711_), .ZN(new_n1712_));
  AOI21_X1  g1334(.A(new_n1422_), .B1(new_n1708_), .B2(new_n1712_), .ZN(new_n1713_));
  NAND2_X1  g1335(.A1(new_n1655_), .A2(new_n794_), .ZN(new_n1714_));
  XNOR2_X1  g1336(.A(new_n682_), .B(new_n665_), .ZN(new_n1715_));
  AOI21_X1  g1337(.A(new_n1427_), .B1(new_n1715_), .B2(new_n680_), .ZN(new_n1716_));
  INV_X1    g1338(.A(new_n1716_), .ZN(new_n1717_));
  AND3_X1   g1339(.A1(new_n1429_), .A2(new_n688_), .A3(new_n1717_), .ZN(new_n1718_));
  AOI21_X1  g1340(.A(new_n1717_), .B1(new_n1429_), .B2(new_n688_), .ZN(new_n1719_));
  NOR3_X1   g1341(.A1(new_n1718_), .A2(new_n1719_), .A3(new_n1434_), .ZN(new_n1720_));
  OAI21_X1  g1342(.A(new_n695_), .B1(new_n1720_), .B2(KEYINPUT58), .ZN(new_n1721_));
  OAI21_X1  g1343(.A(new_n1434_), .B1(new_n1718_), .B2(new_n1719_), .ZN(new_n1722_));
  NAND2_X1  g1344(.A1(new_n1430_), .A2(new_n1716_), .ZN(new_n1723_));
  NAND3_X1  g1345(.A1(new_n1429_), .A2(new_n688_), .A3(new_n1717_), .ZN(new_n1724_));
  NAND3_X1  g1346(.A1(new_n1723_), .A2(new_n675_), .A3(new_n1724_), .ZN(new_n1725_));
  AND3_X1   g1347(.A1(new_n1722_), .A2(new_n1725_), .A3(new_n690_), .ZN(new_n1726_));
  AOI21_X1  g1348(.A(new_n690_), .B1(new_n1722_), .B2(new_n1725_), .ZN(new_n1727_));
  OAI21_X1  g1349(.A(new_n1721_), .B1(new_n1726_), .B2(new_n1727_), .ZN(new_n1728_));
  AOI21_X1  g1350(.A(new_n675_), .B1(new_n1723_), .B2(new_n1724_), .ZN(new_n1729_));
  OAI21_X1  g1351(.A(new_n1698_), .B1(new_n1720_), .B2(new_n1729_), .ZN(new_n1730_));
  INV_X1    g1352(.A(KEYINPUT58), .ZN(new_n1731_));
  AOI21_X1  g1353(.A(new_n774_), .B1(new_n1725_), .B2(new_n1731_), .ZN(new_n1732_));
  NAND3_X1  g1354(.A1(new_n1722_), .A2(new_n1725_), .A3(new_n690_), .ZN(new_n1733_));
  NAND3_X1  g1355(.A1(new_n1730_), .A2(new_n1732_), .A3(new_n1733_), .ZN(new_n1734_));
  AOI21_X1  g1356(.A(new_n1714_), .B1(new_n1728_), .B2(new_n1734_), .ZN(new_n1735_));
  NOR2_X1   g1357(.A1(new_n1713_), .A2(new_n1735_), .ZN(new_n1736_));
  NAND2_X1  g1358(.A1(new_n1728_), .A2(new_n1734_), .ZN(new_n1737_));
  OAI211_X1 g1359(.A(new_n1737_), .B(new_n1389_), .C1(new_n730_), .C2(new_n794_), .ZN(new_n1738_));
  AND2_X1   g1360(.A1(new_n1736_), .A2(new_n1738_), .ZN(new_n1739_));
  NAND4_X1  g1361(.A1(new_n1688_), .A2(new_n1692_), .A3(new_n716_), .A4(new_n1690_), .ZN(new_n1740_));
  INV_X1    g1362(.A(KEYINPUT57), .ZN(new_n1741_));
  NAND2_X1  g1363(.A1(new_n1740_), .A2(new_n1741_), .ZN(new_n1742_));
  NAND3_X1  g1364(.A1(new_n1686_), .A2(new_n1643_), .A3(new_n1687_), .ZN(new_n1743_));
  NAND3_X1  g1365(.A1(new_n1678_), .A2(new_n1683_), .A3(new_n723_), .ZN(new_n1744_));
  NAND3_X1  g1366(.A1(new_n1743_), .A2(new_n1416_), .A3(new_n1744_), .ZN(new_n1745_));
  NAND2_X1  g1367(.A1(new_n1742_), .A2(new_n1745_), .ZN(new_n1746_));
  NOR2_X1   g1368(.A1(new_n1740_), .A2(new_n1741_), .ZN(new_n1747_));
  OAI21_X1  g1369(.A(new_n1389_), .B1(new_n1746_), .B2(new_n1747_), .ZN(new_n1748_));
  INV_X1    g1370(.A(new_n1657_), .ZN(new_n1749_));
  AOI21_X1  g1371(.A(new_n1749_), .B1(new_n1736_), .B2(new_n1738_), .ZN(new_n1750_));
  AOI22_X1  g1372(.A1(new_n1695_), .A2(new_n1739_), .B1(new_n1748_), .B2(new_n1750_), .ZN(G370));
  INV_X1    g1373(.A(KEYINPUT59), .ZN(new_n1752_));
  NAND2_X1  g1374(.A1(new_n635_), .A2(new_n632_), .ZN(new_n1753_));
  OAI21_X1  g1375(.A(new_n1753_), .B1(new_n1110_), .B2(new_n649_), .ZN(new_n1754_));
  OAI211_X1 g1376(.A(new_n1752_), .B(new_n438_), .C1(new_n1104_), .C2(new_n1754_), .ZN(new_n1755_));
  INV_X1    g1377(.A(new_n438_), .ZN(new_n1756_));
  NAND4_X1  g1378(.A1(new_n1098_), .A2(new_n649_), .A3(new_n634_), .A4(new_n650_), .ZN(new_n1757_));
  AOI21_X1  g1379(.A(new_n1756_), .B1(new_n1099_), .B2(new_n1757_), .ZN(new_n1758_));
  OAI21_X1  g1380(.A(KEYINPUT59), .B1(new_n1754_), .B2(new_n438_), .ZN(new_n1759_));
  OAI21_X1  g1381(.A(new_n1755_), .B1(new_n1758_), .B2(new_n1759_), .ZN(new_n1760_));
  NAND2_X1  g1382(.A1(new_n644_), .A2(new_n652_), .ZN(new_n1761_));
  NAND3_X1  g1383(.A1(new_n1093_), .A2(new_n1760_), .A3(new_n1761_), .ZN(new_n1762_));
  NOR2_X1   g1384(.A1(new_n1107_), .A2(new_n652_), .ZN(new_n1763_));
  XOR2_X1   g1385(.A(new_n1763_), .B(new_n439_), .Z(new_n1764_));
  OAI21_X1  g1386(.A(new_n1753_), .B1(new_n636_), .B2(new_n1100_), .ZN(new_n1765_));
  NAND2_X1  g1387(.A1(new_n1765_), .A2(new_n642_), .ZN(new_n1766_));
  NAND4_X1  g1388(.A1(new_n1766_), .A2(new_n641_), .A3(new_n760_), .A4(new_n1761_), .ZN(new_n1767_));
  OAI21_X1  g1389(.A(new_n438_), .B1(new_n1104_), .B2(new_n1754_), .ZN(new_n1768_));
  NAND2_X1  g1390(.A1(new_n1099_), .A2(new_n1756_), .ZN(new_n1769_));
  NAND3_X1  g1391(.A1(new_n1768_), .A2(KEYINPUT59), .A3(new_n1769_), .ZN(new_n1770_));
  NAND3_X1  g1392(.A1(new_n1767_), .A2(new_n1770_), .A3(new_n1755_), .ZN(new_n1771_));
  AND3_X1   g1393(.A1(new_n1762_), .A2(new_n1764_), .A3(new_n1771_), .ZN(new_n1772_));
  AOI21_X1  g1394(.A(new_n1764_), .B1(new_n1762_), .B2(new_n1771_), .ZN(new_n1773_));
  OAI21_X1  g1395(.A(new_n1115_), .B1(new_n1772_), .B2(new_n1773_), .ZN(new_n1774_));
  INV_X1    g1396(.A(new_n1764_), .ZN(new_n1775_));
  AOI21_X1  g1397(.A(new_n1760_), .B1(new_n1093_), .B2(new_n1761_), .ZN(new_n1776_));
  AOI21_X1  g1398(.A(new_n1767_), .B1(new_n1770_), .B2(new_n1755_), .ZN(new_n1777_));
  OAI21_X1  g1399(.A(new_n1775_), .B1(new_n1776_), .B2(new_n1777_), .ZN(new_n1778_));
  NAND3_X1  g1400(.A1(new_n1762_), .A2(new_n1764_), .A3(new_n1771_), .ZN(new_n1779_));
  NAND3_X1  g1401(.A1(new_n1778_), .A2(new_n651_), .A3(new_n1779_), .ZN(new_n1780_));
  NAND3_X1  g1402(.A1(new_n1774_), .A2(new_n1780_), .A3(KEYINPUT60), .ZN(new_n1781_));
  INV_X1    g1403(.A(KEYINPUT60), .ZN(new_n1782_));
  OAI211_X1 g1404(.A(new_n1782_), .B(new_n1115_), .C1(new_n1772_), .C2(new_n1773_), .ZN(new_n1783_));
  AND3_X1   g1405(.A1(new_n1781_), .A2(new_n628_), .A3(new_n1783_), .ZN(new_n1784_));
  AOI21_X1  g1406(.A(new_n628_), .B1(new_n1781_), .B2(new_n1783_), .ZN(new_n1785_));
  NOR2_X1   g1407(.A1(new_n1784_), .A2(new_n1785_), .ZN(new_n1786_));
  AOI21_X1  g1408(.A(new_n629_), .B1(new_n1774_), .B2(new_n1780_), .ZN(new_n1787_));
  OAI21_X1  g1409(.A(new_n636_), .B1(new_n1785_), .B2(new_n1787_), .ZN(new_n1788_));
  INV_X1    g1410(.A(KEYINPUT61), .ZN(new_n1789_));
  AOI22_X1  g1411(.A1(new_n1111_), .A2(new_n1786_), .B1(new_n1788_), .B2(new_n1789_), .ZN(new_n1790_));
  OR2_X1    g1412(.A1(new_n1788_), .A2(new_n1789_), .ZN(new_n1791_));
  AOI21_X1  g1413(.A(new_n752_), .B1(new_n1790_), .B2(new_n1791_), .ZN(new_n1792_));
  OAI21_X1  g1414(.A(new_n1112_), .B1(new_n1784_), .B2(new_n1785_), .ZN(new_n1793_));
  NAND2_X1  g1415(.A1(new_n1781_), .A2(new_n1783_), .ZN(new_n1794_));
  NAND2_X1  g1416(.A1(new_n1794_), .A2(new_n629_), .ZN(new_n1795_));
  INV_X1    g1417(.A(new_n1787_), .ZN(new_n1796_));
  NAND3_X1  g1418(.A1(new_n1795_), .A2(new_n757_), .A3(new_n1796_), .ZN(new_n1797_));
  AND3_X1   g1419(.A1(new_n1793_), .A2(new_n1797_), .A3(new_n752_), .ZN(new_n1798_));
  OAI21_X1  g1420(.A(G4526), .B1(new_n1792_), .B2(new_n1798_), .ZN(new_n1799_));
  XNOR2_X1  g1421(.A(new_n600_), .B(new_n1133_), .ZN(new_n1800_));
  NAND2_X1  g1422(.A1(new_n747_), .A2(new_n748_), .ZN(new_n1801_));
  OAI21_X1  g1423(.A(new_n1801_), .B1(new_n606_), .B2(new_n747_), .ZN(new_n1802_));
  MUX2_X1   g1424(.A(new_n600_), .B(new_n1800_), .S(new_n1802_), .Z(new_n1803_));
  XNOR2_X1  g1425(.A(new_n613_), .B(new_n618_), .ZN(new_n1804_));
  XNOR2_X1  g1426(.A(new_n1803_), .B(new_n1804_), .ZN(new_n1805_));
  INV_X1    g1427(.A(new_n1125_), .ZN(new_n1806_));
  OR2_X1    g1428(.A1(new_n1805_), .A2(new_n1806_), .ZN(new_n1807_));
  NAND2_X1  g1429(.A1(new_n1805_), .A2(new_n1806_), .ZN(new_n1808_));
  NAND3_X1  g1430(.A1(new_n1807_), .A2(new_n1130_), .A3(new_n1808_), .ZN(new_n1809_));
  NAND2_X1  g1431(.A1(new_n1121_), .A2(KEYINPUT63), .ZN(new_n1810_));
  XOR2_X1   g1432(.A(new_n1810_), .B(new_n1804_), .Z(new_n1811_));
  OAI21_X1  g1433(.A(new_n1118_), .B1(new_n604_), .B2(new_n596_), .ZN(new_n1812_));
  OAI21_X1  g1434(.A(new_n1812_), .B1(new_n1121_), .B2(KEYINPUT63), .ZN(new_n1813_));
  XNOR2_X1  g1435(.A(new_n1811_), .B(new_n1813_), .ZN(new_n1814_));
  XNOR2_X1  g1436(.A(new_n1814_), .B(new_n1800_), .ZN(new_n1815_));
  OAI21_X1  g1437(.A(new_n1809_), .B1(new_n1815_), .B2(new_n1130_), .ZN(new_n1816_));
  NAND2_X1  g1438(.A1(new_n1769_), .A2(new_n436_), .ZN(new_n1817_));
  NOR2_X1   g1439(.A1(new_n1099_), .A2(new_n1756_), .ZN(new_n1818_));
  NOR2_X1   g1440(.A1(new_n1817_), .A2(new_n1818_), .ZN(new_n1819_));
  AOI21_X1  g1441(.A(new_n1110_), .B1(new_n1108_), .B2(new_n1753_), .ZN(new_n1820_));
  NOR2_X1   g1442(.A1(new_n1820_), .A2(new_n436_), .ZN(new_n1821_));
  NOR2_X1   g1443(.A1(new_n1819_), .A2(new_n1821_), .ZN(new_n1822_));
  NAND2_X1  g1444(.A1(new_n1093_), .A2(new_n1107_), .ZN(new_n1823_));
  NAND2_X1  g1445(.A1(new_n1766_), .A2(new_n641_), .ZN(new_n1824_));
  NAND2_X1  g1446(.A1(new_n1824_), .A2(new_n1108_), .ZN(new_n1825_));
  NAND3_X1  g1447(.A1(new_n1823_), .A2(new_n651_), .A3(new_n1825_), .ZN(new_n1826_));
  INV_X1    g1448(.A(new_n1826_), .ZN(new_n1827_));
  AOI21_X1  g1449(.A(new_n651_), .B1(new_n1823_), .B2(new_n1825_), .ZN(new_n1828_));
  OAI21_X1  g1450(.A(new_n1822_), .B1(new_n1827_), .B2(new_n1828_), .ZN(new_n1829_));
  INV_X1    g1451(.A(new_n1828_), .ZN(new_n1830_));
  INV_X1    g1452(.A(new_n1822_), .ZN(new_n1831_));
  NAND3_X1  g1453(.A1(new_n1830_), .A2(new_n1826_), .A3(new_n1831_), .ZN(new_n1832_));
  NAND2_X1  g1454(.A1(new_n1829_), .A2(new_n1832_), .ZN(new_n1833_));
  NAND2_X1  g1455(.A1(new_n1833_), .A2(new_n628_), .ZN(new_n1834_));
  NAND3_X1  g1456(.A1(new_n1829_), .A2(new_n1832_), .A3(new_n629_), .ZN(new_n1835_));
  NAND3_X1  g1457(.A1(new_n1834_), .A2(new_n757_), .A3(new_n1835_), .ZN(new_n1836_));
  AND3_X1   g1458(.A1(new_n1834_), .A2(KEYINPUT62), .A3(new_n1835_), .ZN(new_n1837_));
  OAI21_X1  g1459(.A(new_n1112_), .B1(new_n1834_), .B2(KEYINPUT62), .ZN(new_n1838_));
  OAI21_X1  g1460(.A(new_n1836_), .B1(new_n1837_), .B2(new_n1838_), .ZN(new_n1839_));
  AOI21_X1  g1461(.A(G4526), .B1(new_n1839_), .B2(new_n643_), .ZN(new_n1840_));
  OAI211_X1 g1462(.A(new_n752_), .B(new_n1836_), .C1(new_n1837_), .C2(new_n1838_), .ZN(new_n1841_));
  AOI21_X1  g1463(.A(new_n1816_), .B1(new_n1840_), .B2(new_n1841_), .ZN(new_n1842_));
  AOI21_X1  g1464(.A(new_n752_), .B1(new_n1793_), .B2(new_n1797_), .ZN(new_n1843_));
  OAI21_X1  g1465(.A(G4526), .B1(new_n1798_), .B2(new_n1843_), .ZN(new_n1844_));
  NAND2_X1  g1466(.A1(new_n1839_), .A2(new_n643_), .ZN(new_n1845_));
  NAND3_X1  g1467(.A1(new_n1845_), .A2(new_n1102_), .A3(new_n1841_), .ZN(new_n1846_));
  NAND2_X1  g1468(.A1(new_n1844_), .A2(new_n1846_), .ZN(new_n1847_));
  AOI22_X1  g1469(.A1(new_n1799_), .A2(new_n1842_), .B1(new_n1847_), .B2(new_n1816_), .ZN(G399));
endmodule


