//Secret key is'0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_c7552" written by ABC on Wed Nov 16 10:00:29 2022

module locked_c7552 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G5, G9, G12, G15, G18, G23, G26, G29,
    G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59,
    G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77,
    G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97,
    G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121,
    G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151,
    G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163,
    G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175,
    G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187,
    G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199,
    G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211,
    G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223,
    G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235,
    G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469,
    G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230,
    G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717,
    G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410,
    G4415, G4420, G4427, G4432, G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G5, G9, G12, G15, G18, G23,
    G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57,
    G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75,
    G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89,
    G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115,
    G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147,
    G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161,
    G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173,
    G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185,
    G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197,
    G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209,
    G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221,
    G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233,
    G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459,
    G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218,
    G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705,
    G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400,
    G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_n484_, new_n491_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1256_, new_n1258_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1446_, new_n1448_, new_n1449_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1470_, new_n1471_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1482_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1511_,
    new_n1512_, new_n1513_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1540_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_;
  BUF_X1    g0000(.A(G1), .Z(G2));
  BUF_X1    g0001(.A(G1), .Z(G3));
  XOR2_X1   g0002(.A(KEYINPUT0), .B(G1459), .Z(G450));
  BUF_X1    g0003(.A(G1469), .Z(G448));
  BUF_X1    g0004(.A(G1480), .Z(G444));
  BUF_X1    g0005(.A(G1486), .Z(G442));
  BUF_X1    g0006(.A(G1492), .Z(G440));
  BUF_X1    g0007(.A(G1496), .Z(G438));
  BUF_X1    g0008(.A(G2208), .Z(G496));
  BUF_X1    g0009(.A(G2218), .Z(G494));
  BUF_X1    g0010(.A(G2224), .Z(G492));
  BUF_X1    g0011(.A(G2230), .Z(G490));
  BUF_X1    g0012(.A(G2236), .Z(G488));
  BUF_X1    g0013(.A(G2239), .Z(G486));
  BUF_X1    g0014(.A(G2247), .Z(G484));
  BUF_X1    g0015(.A(G2253), .Z(G482));
  BUF_X1    g0016(.A(G2256), .Z(G480));
  BUF_X1    g0017(.A(G3698), .Z(G560));
  BUF_X1    g0018(.A(G3701), .Z(G542));
  BUF_X1    g0019(.A(G3705), .Z(G558));
  BUF_X1    g0020(.A(G3711), .Z(G556));
  BUF_X1    g0021(.A(G3717), .Z(G554));
  BUF_X1    g0022(.A(G3723), .Z(G552));
  BUF_X1    g0023(.A(G3729), .Z(G550));
  BUF_X1    g0024(.A(G3737), .Z(G548));
  BUF_X1    g0025(.A(G3743), .Z(G546));
  BUF_X1    g0026(.A(G3749), .Z(G544));
  BUF_X1    g0027(.A(G4393), .Z(G540));
  BUF_X1    g0028(.A(G4400), .Z(G538));
  BUF_X1    g0029(.A(G4405), .Z(G536));
  BUF_X1    g0030(.A(G4410), .Z(G534));
  BUF_X1    g0031(.A(G4415), .Z(G532));
  BUF_X1    g0032(.A(G4420), .Z(G530));
  BUF_X1    g0033(.A(G4427), .Z(G528));
  XNOR2_X1  g0034(.A(KEYINPUT1), .B(G4432), .ZN(G526));
  BUF_X1    g0035(.A(G4437), .Z(G524));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G15), .ZN(G279));
  BUF_X1    g0037(.A(G1462), .Z(G436));
  BUF_X1    g0038(.A(G2211), .Z(G478));
  BUF_X1    g0039(.A(G4394), .Z(G522));
  OR2_X1    g0040(.A1(G5), .A2(G57), .ZN(G402));
  NAND4_X1  g0041(.A1(G150), .A2(G184), .A3(G228), .A4(G240), .ZN(new_n484_));
  XOR2_X1   g0042(.A(new_n484_), .B(KEYINPUT3), .Z(G404));
  NAND4_X1  g0043(.A1(G152), .A2(G210), .A3(G218), .A4(G230), .ZN(G406));
  NAND4_X1  g0044(.A1(G182), .A2(G183), .A3(G185), .A4(G186), .ZN(G408));
  NAND4_X1  g0045(.A1(G162), .A2(G172), .A3(G188), .A4(G199), .ZN(G410));
  BUF_X1    g0046(.A(G1), .Z(G432));
  BUF_X1    g0047(.A(G106), .Z(G446));
  INV_X1    g0048(.A(G5), .ZN(new_n491_));
  NAND2_X1  g0049(.A1(new_n491_), .A2(G1197), .ZN(G284));
  INV_X1    g0050(.A(G15), .ZN(G286));
  NAND2_X1  g0051(.A1(new_n491_), .A2(G1197), .ZN(G289));
  NAND3_X1  g0052(.A1(new_n491_), .A2(G133), .A3(G134), .ZN(G292));
  INV_X1    g0053(.A(G15), .ZN(G341));
  NAND3_X1  g0054(.A1(new_n491_), .A2(G133), .A3(G134), .ZN(G281));
  BUF_X1    g0055(.A(G1), .Z(G453));
  AND2_X1   g0056(.A1(G1), .A2(G163), .ZN(G278));
  INV_X1    g0057(.A(G41), .ZN(new_n500_));
  NOR3_X1   g0058(.A1(new_n500_), .A2(G18), .A3(G3701), .ZN(new_n501_));
  INV_X1    g0059(.A(G3701), .ZN(new_n502_));
  NOR3_X1   g0060(.A1(new_n502_), .A2(G18), .A3(G41), .ZN(new_n503_));
  NOR2_X1   g0061(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g0062(.A(G4526), .ZN(new_n505_));
  XNOR2_X1  g0063(.A(new_n504_), .B(new_n505_), .ZN(G373));
  INV_X1    g0064(.A(G18), .ZN(new_n507_));
  AND2_X1   g0065(.A1(new_n507_), .A2(G50), .ZN(new_n508_));
  AOI21_X1  g0066(.A(new_n508_), .B1(G18), .B2(G220), .ZN(new_n509_));
  NOR2_X1   g0067(.A1(new_n509_), .A2(G4432), .ZN(new_n510_));
  INV_X1    g0068(.A(G4427), .ZN(new_n511_));
  INV_X1    g0069(.A(G32), .ZN(new_n512_));
  NOR2_X1   g0070(.A1(new_n512_), .A2(G18), .ZN(new_n513_));
  AND2_X1   g0071(.A1(G18), .A2(G221), .ZN(new_n514_));
  OAI21_X1  g0072(.A(new_n511_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g0073(.A(new_n515_), .B(KEYINPUT30), .ZN(new_n516_));
  NAND2_X1  g0074(.A1(new_n509_), .A2(G4432), .ZN(new_n517_));
  AOI21_X1  g0075(.A(new_n510_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g0076(.A(new_n517_), .ZN(new_n519_));
  NOR2_X1   g0077(.A1(new_n519_), .A2(new_n510_), .ZN(new_n520_));
  AOI21_X1  g0078(.A(new_n513_), .B1(G18), .B2(G221), .ZN(new_n521_));
  NAND2_X1  g0079(.A1(new_n521_), .A2(G4427), .ZN(new_n522_));
  AND2_X1   g0080(.A1(new_n522_), .A2(new_n515_), .ZN(new_n523_));
  NAND2_X1  g0081(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g0082(.A1(new_n507_), .A2(G35), .ZN(new_n525_));
  INV_X1    g0083(.A(G222), .ZN(new_n526_));
  OAI21_X1  g0084(.A(new_n525_), .B1(new_n507_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g0085(.A(G4420), .ZN(new_n528_));
  NAND2_X1  g0086(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g0087(.A(new_n518_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g0088(.A(G66), .ZN(new_n531_));
  NOR2_X1   g0089(.A1(new_n531_), .A2(G18), .ZN(new_n532_));
  AOI21_X1  g0090(.A(new_n532_), .B1(G18), .B2(G219), .ZN(new_n533_));
  NAND2_X1  g0091(.A1(new_n533_), .A2(G4437), .ZN(new_n534_));
  NAND2_X1  g0092(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  OR2_X1    g0093(.A1(new_n533_), .A2(G4437), .ZN(new_n536_));
  NAND2_X1  g0094(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g0095(.A1(G18), .A2(G223), .ZN(new_n538_));
  INV_X1    g0096(.A(G47), .ZN(new_n539_));
  OAI21_X1  g0097(.A(new_n538_), .B1(new_n539_), .B2(G18), .ZN(new_n540_));
  INV_X1    g0098(.A(G4415), .ZN(new_n541_));
  OR2_X1    g0099(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g0100(.A1(new_n540_), .A2(new_n541_), .ZN(new_n543_));
  NAND2_X1  g0101(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g0102(.A1(G18), .A2(G225), .ZN(new_n545_));
  INV_X1    g0103(.A(G94), .ZN(new_n546_));
  OAI21_X1  g0104(.A(new_n545_), .B1(new_n546_), .B2(G18), .ZN(new_n547_));
  INV_X1    g0105(.A(G4405), .ZN(new_n548_));
  NAND2_X1  g0106(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g0107(.A1(new_n507_), .A2(G118), .ZN(new_n550_));
  INV_X1    g0108(.A(G217), .ZN(new_n551_));
  OAI21_X1  g0109(.A(new_n550_), .B1(new_n507_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g0110(.A(new_n552_), .ZN(new_n553_));
  OR2_X1    g0111(.A1(new_n553_), .A2(G4394), .ZN(new_n554_));
  NAND2_X1  g0112(.A1(G18), .A2(G226), .ZN(new_n555_));
  INV_X1    g0113(.A(G97), .ZN(new_n556_));
  OAI21_X1  g0114(.A(new_n555_), .B1(new_n556_), .B2(G18), .ZN(new_n557_));
  INV_X1    g0115(.A(G4400), .ZN(new_n558_));
  OR2_X1    g0116(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g0117(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g0118(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OR2_X1    g0119(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g0120(.A(new_n547_), .B(G4405), .ZN(new_n563_));
  INV_X1    g0121(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g0122(.A(new_n549_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g0123(.A1(new_n507_), .A2(G121), .ZN(new_n566_));
  INV_X1    g0124(.A(G224), .ZN(new_n567_));
  OAI21_X1  g0125(.A(new_n566_), .B1(new_n507_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g0126(.A(new_n568_), .B(G4410), .ZN(new_n569_));
  NAND2_X1  g0127(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g0128(.A(new_n560_), .B(KEYINPUT26), .ZN(new_n571_));
  NAND3_X1  g0129(.A1(new_n571_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n572_));
  INV_X1    g0130(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g0131(.A1(new_n573_), .A2(KEYINPUT27), .ZN(new_n574_));
  AOI21_X1  g0132(.A(new_n544_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g0133(.A(new_n543_), .B(KEYINPUT25), .Z(new_n576_));
  XNOR2_X1  g0134(.A(new_n544_), .B(KEYINPUT28), .ZN(new_n577_));
  INV_X1    g0135(.A(G4410), .ZN(new_n578_));
  NAND2_X1  g0136(.A1(new_n568_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g0137(.A1(new_n572_), .A2(new_n544_), .ZN(new_n580_));
  OAI221_X1 g0138(.A(new_n576_), .B1(new_n577_), .B2(new_n579_), .C1(new_n580_), .C2(KEYINPUT27), .ZN(new_n581_));
  NOR2_X1   g0139(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g0140(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g0141(.A(new_n520_), .ZN(new_n584_));
  XNOR2_X1  g0142(.A(KEYINPUT19), .B(G4420), .ZN(new_n585_));
  XOR2_X1   g0143(.A(new_n527_), .B(new_n585_), .Z(new_n586_));
  NAND2_X1  g0144(.A1(new_n536_), .A2(new_n534_), .ZN(new_n587_));
  NOR3_X1   g0145(.A1(new_n584_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g0146(.A(new_n523_), .B(KEYINPUT18), .ZN(new_n589_));
  AND2_X1   g0147(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g0148(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g0149(.A(new_n591_), .B(KEYINPUT29), .ZN(new_n592_));
  NAND2_X1  g0150(.A1(new_n507_), .A2(G100), .ZN(new_n593_));
  NAND2_X1  g0151(.A1(G18), .A2(G231), .ZN(new_n594_));
  AND2_X1   g0152(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OR2_X1    g0153(.A1(new_n595_), .A2(G3749), .ZN(new_n596_));
  INV_X1    g0154(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g0155(.A1(new_n507_), .A2(G124), .ZN(new_n598_));
  NAND2_X1  g0156(.A1(G18), .A2(G232), .ZN(new_n599_));
  AND2_X1   g0157(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OR2_X1    g0158(.A1(new_n600_), .A2(G3743), .ZN(new_n601_));
  NAND2_X1  g0159(.A1(new_n600_), .A2(G3743), .ZN(new_n602_));
  AND2_X1   g0160(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g0161(.A(new_n603_), .B(KEYINPUT16), .ZN(new_n604_));
  AND2_X1   g0162(.A1(new_n507_), .A2(G127), .ZN(new_n605_));
  AOI21_X1  g0163(.A(new_n605_), .B1(G18), .B2(G233), .ZN(new_n606_));
  NOR2_X1   g0164(.A1(new_n606_), .A2(G3737), .ZN(new_n607_));
  INV_X1    g0165(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g0166(.A1(new_n606_), .A2(G3737), .ZN(new_n609_));
  AND2_X1   g0167(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g0168(.A1(new_n507_), .A2(G130), .ZN(new_n611_));
  NAND2_X1  g0169(.A1(G18), .A2(G234), .ZN(new_n612_));
  AND2_X1   g0170(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OR2_X1    g0171(.A1(new_n613_), .A2(G3729), .ZN(new_n614_));
  INV_X1    g0172(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g0173(.A1(new_n604_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g0174(.A(new_n601_), .B(KEYINPUT17), .ZN(new_n617_));
  AOI21_X1  g0175(.A(new_n617_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n618_));
  NAND2_X1  g0176(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g0177(.A1(new_n595_), .A2(G3749), .ZN(new_n620_));
  AOI21_X1  g0178(.A(new_n597_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g0179(.A(new_n621_), .ZN(new_n622_));
  AND2_X1   g0180(.A1(G18), .A2(G235), .ZN(new_n623_));
  AOI21_X1  g0181(.A(new_n623_), .B1(new_n507_), .B2(G103), .ZN(new_n624_));
  NOR2_X1   g0182(.A1(new_n624_), .A2(G3723), .ZN(new_n625_));
  NAND2_X1  g0183(.A1(new_n507_), .A2(G23), .ZN(new_n626_));
  INV_X1    g0184(.A(G236), .ZN(new_n627_));
  OAI21_X1  g0185(.A(new_n626_), .B1(new_n507_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g0186(.A(KEYINPUT11), .ZN(new_n629_));
  INV_X1    g0187(.A(G3717), .ZN(new_n630_));
  NOR2_X1   g0188(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OR2_X1    g0189(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g0190(.A1(KEYINPUT11), .A2(G3717), .ZN(new_n633_));
  OAI21_X1  g0191(.A(new_n628_), .B1(new_n633_), .B2(new_n631_), .ZN(new_n634_));
  NAND2_X1  g0192(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g0193(.A1(new_n507_), .A2(G26), .ZN(new_n636_));
  INV_X1    g0194(.A(G237), .ZN(new_n637_));
  OAI21_X1  g0195(.A(new_n636_), .B1(new_n507_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g0196(.A1(new_n638_), .A2(G3711), .ZN(new_n639_));
  INV_X1    g0197(.A(KEYINPUT12), .ZN(new_n640_));
  INV_X1    g0198(.A(G3711), .ZN(new_n641_));
  OAI211_X1 g0199(.A(new_n636_), .B(new_n641_), .C1(new_n507_), .C2(new_n637_), .ZN(new_n642_));
  NAND3_X1  g0200(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g0201(.A1(new_n638_), .A2(KEYINPUT12), .A3(G3711), .ZN(new_n644_));
  NAND2_X1  g0202(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g0203(.A(KEYINPUT13), .B1(G18), .B2(G238), .ZN(new_n646_));
  NAND2_X1  g0204(.A1(new_n507_), .A2(G29), .ZN(new_n647_));
  NAND2_X1  g0205(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g0206(.A(G3705), .ZN(new_n649_));
  NAND3_X1  g0207(.A1(KEYINPUT13), .A2(G18), .A3(G238), .ZN(new_n650_));
  NAND3_X1  g0208(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g0209(.A(new_n651_), .B(KEYINPUT15), .ZN(new_n652_));
  XOR2_X1   g0210(.A(KEYINPUT14), .B(G3705), .Z(new_n653_));
  INV_X1    g0211(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g0212(.A1(new_n648_), .A2(new_n650_), .ZN(new_n655_));
  NAND2_X1  g0213(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g0214(.A1(new_n656_), .A2(new_n501_), .A3(new_n651_), .ZN(new_n657_));
  AOI21_X1  g0215(.A(new_n645_), .B1(new_n652_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g0216(.A1(new_n638_), .A2(new_n641_), .ZN(new_n659_));
  INV_X1    g0217(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g0218(.A(new_n635_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0219(.A1(new_n628_), .A2(new_n630_), .ZN(new_n662_));
  NAND2_X1  g0220(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g0221(.A1(new_n624_), .A2(G3723), .ZN(new_n664_));
  AOI21_X1  g0222(.A(new_n625_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g0223(.A1(new_n656_), .A2(new_n504_), .A3(new_n651_), .ZN(new_n666_));
  NOR2_X1   g0224(.A1(new_n666_), .A2(new_n505_), .ZN(new_n667_));
  INV_X1    g0225(.A(new_n645_), .ZN(new_n668_));
  INV_X1    g0226(.A(new_n664_), .ZN(new_n669_));
  NOR2_X1   g0227(.A1(new_n669_), .A2(new_n625_), .ZN(new_n670_));
  NAND4_X1  g0228(.A1(new_n667_), .A2(new_n668_), .A3(new_n670_), .A4(new_n635_), .ZN(new_n671_));
  NAND2_X1  g0229(.A1(new_n665_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g0230(.A1(new_n596_), .A2(new_n620_), .ZN(new_n673_));
  NAND2_X1  g0231(.A1(new_n613_), .A2(G3729), .ZN(new_n674_));
  NAND2_X1  g0232(.A1(new_n614_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g0233(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  AND3_X1   g0234(.A1(new_n604_), .A2(new_n610_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g0235(.A(new_n622_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g0236(.A1(new_n553_), .A2(G4394), .ZN(new_n679_));
  NAND2_X1  g0237(.A1(new_n554_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g0238(.A1(new_n680_), .A2(new_n561_), .ZN(new_n681_));
  NAND3_X1  g0239(.A1(new_n681_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n682_));
  NOR3_X1   g0240(.A1(new_n678_), .A2(new_n682_), .A3(new_n544_), .ZN(new_n683_));
  AOI211_X1 g0241(.A(new_n537_), .B(new_n592_), .C1(new_n590_), .C2(new_n683_), .ZN(new_n684_));
  AND2_X1   g0242(.A1(G9), .A2(G12), .ZN(new_n685_));
  INV_X1    g0243(.A(G154), .ZN(new_n686_));
  AOI21_X1  g0244(.A(new_n685_), .B1(G18), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g0245(.A(G2253), .ZN(new_n688_));
  NAND2_X1  g0246(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g0247(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g0248(.A1(new_n687_), .A2(new_n688_), .ZN(new_n691_));
  NOR2_X1   g0249(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g0250(.A(new_n692_), .B(KEYINPUT5), .Z(new_n693_));
  OR2_X1    g0251(.A1(new_n507_), .A2(G156), .ZN(new_n694_));
  NAND2_X1  g0252(.A1(G9), .A2(G12), .ZN(new_n695_));
  AND2_X1   g0253(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g0254(.A(G2239), .ZN(new_n697_));
  NAND2_X1  g0255(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g0256(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g0257(.A1(new_n694_), .A2(new_n695_), .ZN(new_n700_));
  NAND2_X1  g0258(.A1(new_n700_), .A2(G2239), .ZN(new_n701_));
  INV_X1    g0259(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g0260(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g0261(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g0262(.A(new_n695_), .B1(new_n507_), .B2(G153), .ZN(new_n705_));
  XNOR2_X1  g0263(.A(new_n705_), .B(KEYINPUT7), .ZN(new_n706_));
  NOR2_X1   g0264(.A1(new_n706_), .A2(G2256), .ZN(new_n707_));
  INV_X1    g0265(.A(new_n707_), .ZN(new_n708_));
  NAND2_X1  g0266(.A1(new_n706_), .A2(G2256), .ZN(new_n709_));
  NAND2_X1  g0267(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g0268(.A(new_n695_), .B1(new_n507_), .B2(G155), .ZN(new_n711_));
  INV_X1    g0269(.A(KEYINPUT6), .ZN(new_n712_));
  XNOR2_X1  g0270(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND2_X1  g0271(.A1(new_n713_), .A2(G2247), .ZN(new_n714_));
  OR2_X1    g0272(.A1(new_n711_), .A2(G2247), .ZN(new_n715_));
  NAND2_X1  g0273(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NOR4_X1   g0274(.A1(new_n693_), .A2(new_n704_), .A3(new_n710_), .A4(new_n716_), .ZN(new_n717_));
  INV_X1    g0275(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g0276(.A1(new_n507_), .A2(G144), .ZN(new_n719_));
  NAND2_X1  g0277(.A1(G18), .A2(G159), .ZN(new_n720_));
  AOI21_X1  g0278(.A(G2224), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g0279(.A(new_n721_), .ZN(new_n722_));
  INV_X1    g0280(.A(G144), .ZN(new_n723_));
  OAI211_X1 g0281(.A(new_n720_), .B(G2224), .C1(G18), .C2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g0282(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g0283(.A1(G18), .A2(G158), .ZN(new_n726_));
  INV_X1    g0284(.A(G2230), .ZN(new_n727_));
  INV_X1    g0285(.A(G135), .ZN(new_n728_));
  OAI211_X1 g0286(.A(new_n726_), .B(new_n727_), .C1(G18), .C2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g0287(.A1(new_n729_), .A2(KEYINPUT9), .ZN(new_n730_));
  NAND2_X1  g0288(.A1(new_n507_), .A2(G135), .ZN(new_n731_));
  INV_X1    g0289(.A(KEYINPUT9), .ZN(new_n732_));
  NAND4_X1  g0290(.A1(new_n731_), .A2(new_n732_), .A3(new_n727_), .A4(new_n726_), .ZN(new_n733_));
  AND2_X1   g0291(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g0292(.A1(new_n731_), .A2(new_n726_), .ZN(new_n735_));
  NAND2_X1  g0293(.A1(new_n735_), .A2(KEYINPUT8), .ZN(new_n736_));
  INV_X1    g0294(.A(KEYINPUT8), .ZN(new_n737_));
  OAI211_X1 g0295(.A(new_n726_), .B(new_n737_), .C1(G18), .C2(new_n728_), .ZN(new_n738_));
  NAND3_X1  g0296(.A1(new_n736_), .A2(G2230), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g0297(.A(new_n725_), .B1(new_n734_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g0298(.A(G2211), .ZN(new_n741_));
  NAND2_X1  g0299(.A1(G18), .A2(G151), .ZN(new_n742_));
  INV_X1    g0300(.A(new_n742_), .ZN(new_n743_));
  INV_X1    g0301(.A(G147), .ZN(new_n744_));
  OAI21_X1  g0302(.A(KEYINPUT10), .B1(new_n744_), .B2(G18), .ZN(new_n745_));
  INV_X1    g0303(.A(KEYINPUT10), .ZN(new_n746_));
  NAND3_X1  g0304(.A1(new_n746_), .A2(new_n507_), .A3(G147), .ZN(new_n747_));
  AOI211_X1 g0305(.A(new_n741_), .B(new_n743_), .C1(new_n745_), .C2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g0306(.A1(new_n745_), .A2(new_n747_), .ZN(new_n749_));
  AOI21_X1  g0307(.A(G2211), .B1(new_n749_), .B2(new_n742_), .ZN(new_n750_));
  NAND2_X1  g0308(.A1(G18), .A2(G160), .ZN(new_n751_));
  INV_X1    g0309(.A(G138), .ZN(new_n752_));
  OAI21_X1  g0310(.A(new_n751_), .B1(new_n752_), .B2(G18), .ZN(new_n753_));
  INV_X1    g0311(.A(G2218), .ZN(new_n754_));
  NAND2_X1  g0312(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g0313(.A1(new_n507_), .A2(G138), .ZN(new_n756_));
  NAND3_X1  g0314(.A1(new_n756_), .A2(G2218), .A3(new_n751_), .ZN(new_n757_));
  NAND2_X1  g0315(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g0316(.A1(new_n748_), .A2(new_n750_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g0317(.A1(new_n740_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g0318(.A(new_n695_), .B1(new_n507_), .B2(G157), .ZN(new_n761_));
  INV_X1    g0319(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g0320(.A(G2236), .ZN(new_n763_));
  NAND2_X1  g0321(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g0322(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g0323(.A1(new_n762_), .A2(new_n763_), .ZN(new_n766_));
  NOR2_X1   g0324(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g0325(.A(new_n767_), .ZN(new_n768_));
  NOR2_X1   g0326(.A1(new_n760_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g0327(.A(new_n769_), .ZN(new_n770_));
  NOR3_X1   g0328(.A1(new_n684_), .A2(new_n718_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g0329(.A(G214), .ZN(new_n772_));
  AOI21_X1  g0330(.A(new_n685_), .B1(G18), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g0331(.A(G1480), .ZN(new_n774_));
  NAND2_X1  g0332(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g0333(.A(new_n775_), .ZN(new_n776_));
  NOR2_X1   g0334(.A1(new_n773_), .A2(new_n774_), .ZN(new_n777_));
  NOR2_X1   g0335(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g0336(.A(new_n778_), .ZN(new_n779_));
  OAI21_X1  g0337(.A(new_n695_), .B1(new_n507_), .B2(G215), .ZN(new_n780_));
  INV_X1    g0338(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g0339(.A(G106), .ZN(new_n782_));
  AND2_X1   g0340(.A1(new_n782_), .A2(KEYINPUT4), .ZN(new_n783_));
  NOR2_X1   g0341(.A1(new_n782_), .A2(KEYINPUT4), .ZN(new_n784_));
  OAI21_X1  g0342(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g0343(.A(new_n780_), .B1(KEYINPUT4), .B2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g0344(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g0345(.A(new_n787_), .ZN(new_n788_));
  NOR2_X1   g0346(.A1(new_n779_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g0347(.A(new_n695_), .B1(new_n507_), .B2(G216), .ZN(new_n790_));
  INV_X1    g0348(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g0349(.A(G1469), .ZN(new_n792_));
  NAND2_X1  g0350(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g0351(.A1(new_n790_), .A2(G1469), .ZN(new_n794_));
  NAND2_X1  g0352(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g0353(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g0354(.A(G209), .ZN(new_n797_));
  AOI21_X1  g0355(.A(new_n685_), .B1(G18), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g0356(.A(G1462), .ZN(new_n799_));
  NAND2_X1  g0357(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g0358(.A(new_n800_), .ZN(new_n801_));
  NOR2_X1   g0359(.A1(new_n798_), .A2(new_n799_), .ZN(new_n802_));
  NOR2_X1   g0360(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g0361(.A1(new_n789_), .A2(new_n796_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g0362(.A(G213), .ZN(new_n805_));
  AOI21_X1  g0363(.A(new_n685_), .B1(G18), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g0364(.A(G1486), .ZN(new_n807_));
  NAND2_X1  g0365(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g0366(.A(new_n808_), .ZN(new_n809_));
  NOR2_X1   g0367(.A1(new_n806_), .A2(new_n807_), .ZN(new_n810_));
  NOR2_X1   g0368(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g0369(.A(new_n811_), .ZN(new_n812_));
  NOR2_X1   g0370(.A1(new_n804_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g0371(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g0372(.A1(G1496), .A2(G4528), .ZN(new_n815_));
  NAND2_X1  g0373(.A1(new_n815_), .A2(G38), .ZN(new_n816_));
  INV_X1    g0374(.A(G38), .ZN(new_n817_));
  NAND3_X1  g0375(.A1(new_n817_), .A2(G1496), .A3(G4528), .ZN(new_n818_));
  NAND2_X1  g0376(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g0377(.A1(G1492), .A2(G4528), .ZN(new_n820_));
  NAND2_X1  g0378(.A1(new_n820_), .A2(G38), .ZN(new_n821_));
  NAND3_X1  g0379(.A1(new_n817_), .A2(G1492), .A3(G4528), .ZN(new_n822_));
  NAND2_X1  g0380(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OR2_X1    g0381(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g0382(.A1(new_n814_), .A2(new_n824_), .ZN(new_n825_));
  AND2_X1   g0383(.A1(new_n771_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g0384(.A1(new_n713_), .A2(G2247), .ZN(new_n827_));
  NOR2_X1   g0385(.A1(new_n827_), .A2(new_n690_), .ZN(new_n828_));
  NAND3_X1  g0386(.A1(new_n714_), .A2(new_n699_), .A3(new_n715_), .ZN(new_n829_));
  AOI21_X1  g0387(.A(new_n691_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g0388(.A(new_n707_), .B1(new_n830_), .B2(new_n709_), .ZN(new_n831_));
  AOI211_X1 g0389(.A(KEYINPUT20), .B(G2218), .C1(new_n756_), .C2(new_n751_), .ZN(new_n832_));
  INV_X1    g0390(.A(KEYINPUT20), .ZN(new_n833_));
  AOI21_X1  g0391(.A(new_n833_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n834_));
  NOR2_X1   g0392(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g0393(.A(new_n721_), .B1(new_n835_), .B2(new_n724_), .ZN(new_n836_));
  INV_X1    g0394(.A(new_n757_), .ZN(new_n837_));
  AOI21_X1  g0395(.A(G2218), .B1(new_n756_), .B2(new_n751_), .ZN(new_n838_));
  NOR2_X1   g0396(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g0397(.A(new_n724_), .ZN(new_n840_));
  NOR2_X1   g0398(.A1(new_n840_), .A2(new_n721_), .ZN(new_n841_));
  NAND3_X1  g0399(.A1(new_n839_), .A2(new_n750_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g0400(.A1(new_n836_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g0401(.A(new_n738_), .ZN(new_n844_));
  AOI21_X1  g0402(.A(new_n737_), .B1(new_n731_), .B2(new_n726_), .ZN(new_n845_));
  NOR3_X1   g0403(.A1(new_n844_), .A2(new_n845_), .A3(new_n727_), .ZN(new_n846_));
  NAND2_X1  g0404(.A1(new_n730_), .A2(new_n733_), .ZN(new_n847_));
  NOR2_X1   g0405(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g0406(.A1(new_n848_), .A2(new_n766_), .ZN(new_n849_));
  AOI21_X1  g0407(.A(new_n765_), .B1(new_n843_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g0408(.A(KEYINPUT21), .ZN(new_n851_));
  OR2_X1    g0409(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g0410(.A1(new_n736_), .A2(new_n738_), .ZN(new_n853_));
  NOR2_X1   g0411(.A1(new_n853_), .A2(G2230), .ZN(new_n854_));
  AOI22_X1  g0412(.A1(new_n850_), .A2(new_n851_), .B1(new_n767_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g0413(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g0414(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g0415(.A(new_n831_), .B1(new_n857_), .B2(new_n718_), .ZN(new_n858_));
  NAND2_X1  g0416(.A1(new_n858_), .A2(new_n825_), .ZN(new_n859_));
  XOR2_X1   g0417(.A(new_n859_), .B(KEYINPUT22), .Z(new_n860_));
  OAI21_X1  g0418(.A(G38), .B1(new_n815_), .B2(new_n820_), .ZN(new_n861_));
  XNOR2_X1  g0419(.A(new_n861_), .B(KEYINPUT23), .ZN(new_n862_));
  NAND2_X1  g0420(.A1(new_n796_), .A2(new_n801_), .ZN(new_n863_));
  INV_X1    g0421(.A(KEYINPUT24), .ZN(new_n864_));
  NAND2_X1  g0422(.A1(new_n793_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g0423(.A1(new_n791_), .A2(KEYINPUT24), .A3(new_n792_), .ZN(new_n866_));
  NAND2_X1  g0424(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g0425(.A1(new_n863_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g0426(.A1(new_n868_), .A2(new_n811_), .A3(new_n778_), .A4(new_n787_), .ZN(new_n869_));
  INV_X1    g0427(.A(new_n810_), .ZN(new_n870_));
  NAND2_X1  g0428(.A1(new_n781_), .A2(new_n782_), .ZN(new_n871_));
  AOI21_X1  g0429(.A(new_n777_), .B1(new_n775_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g0430(.A(new_n870_), .B1(new_n872_), .B2(new_n809_), .ZN(new_n873_));
  NAND2_X1  g0431(.A1(new_n869_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g0432(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g0433(.A(new_n862_), .B1(new_n875_), .B2(new_n824_), .ZN(new_n876_));
  OR3_X1    g0434(.A1(new_n826_), .A2(new_n860_), .A3(new_n876_), .ZN(G246));
  OAI21_X1  g0435(.A(new_n695_), .B1(new_n507_), .B2(G173), .ZN(new_n878_));
  XNOR2_X1  g0436(.A(new_n878_), .B(KEYINPUT38), .ZN(new_n879_));
  NOR2_X1   g0437(.A1(G18), .A2(G110), .ZN(new_n880_));
  AOI21_X1  g0438(.A(new_n880_), .B1(G18), .B2(G2256), .ZN(new_n881_));
  NAND2_X1  g0439(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g0440(.A(new_n882_), .B(KEYINPUT47), .ZN(new_n883_));
  XOR2_X1   g0441(.A(new_n879_), .B(new_n881_), .Z(new_n884_));
  OR2_X1    g0442(.A1(new_n507_), .A2(G175), .ZN(new_n885_));
  NAND2_X1  g0443(.A1(new_n885_), .A2(new_n695_), .ZN(new_n886_));
  NOR2_X1   g0444(.A1(G18), .A2(G86), .ZN(new_n887_));
  AOI21_X1  g0445(.A(new_n887_), .B1(G18), .B2(G2247), .ZN(new_n888_));
  INV_X1    g0446(.A(new_n888_), .ZN(new_n889_));
  NOR2_X1   g0447(.A1(G18), .A2(G109), .ZN(new_n890_));
  AOI21_X1  g0448(.A(new_n890_), .B1(G18), .B2(G2253), .ZN(new_n891_));
  INV_X1    g0449(.A(new_n891_), .ZN(new_n892_));
  OAI21_X1  g0450(.A(new_n695_), .B1(new_n507_), .B2(G174), .ZN(new_n893_));
  OAI22_X1  g0451(.A1(new_n886_), .A2(new_n889_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g0452(.A1(new_n892_), .A2(new_n893_), .ZN(new_n895_));
  NAND3_X1  g0453(.A1(new_n884_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g0454(.A(new_n894_), .ZN(new_n897_));
  NAND2_X1  g0455(.A1(new_n889_), .A2(new_n886_), .ZN(new_n898_));
  NAND4_X1  g0456(.A1(new_n884_), .A2(new_n897_), .A3(new_n898_), .A4(new_n895_), .ZN(new_n899_));
  OAI21_X1  g0457(.A(new_n695_), .B1(new_n507_), .B2(G176), .ZN(new_n900_));
  INV_X1    g0458(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g0459(.A1(G18), .A2(G63), .ZN(new_n902_));
  AOI21_X1  g0460(.A(new_n902_), .B1(G18), .B2(G2239), .ZN(new_n903_));
  NAND2_X1  g0461(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g0462(.A(new_n883_), .B(new_n896_), .C1(new_n899_), .C2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g0463(.A(new_n695_), .B1(new_n507_), .B2(G177), .ZN(new_n906_));
  NAND2_X1  g0464(.A1(G18), .A2(G2236), .ZN(new_n907_));
  OAI21_X1  g0465(.A(new_n907_), .B1(G18), .B2(G64), .ZN(new_n908_));
  OR2_X1    g0466(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g0467(.A(new_n906_), .B(new_n908_), .ZN(new_n910_));
  XOR2_X1   g0468(.A(new_n910_), .B(KEYINPUT37), .Z(new_n911_));
  INV_X1    g0469(.A(new_n911_), .ZN(new_n912_));
  INV_X1    g0470(.A(new_n756_), .ZN(new_n913_));
  AOI21_X1  g0471(.A(new_n913_), .B1(G18), .B2(G180), .ZN(new_n914_));
  INV_X1    g0472(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g0473(.A1(G18), .A2(G83), .ZN(new_n916_));
  AOI21_X1  g0474(.A(new_n916_), .B1(G18), .B2(G2218), .ZN(new_n917_));
  INV_X1    g0475(.A(new_n719_), .ZN(new_n918_));
  AOI21_X1  g0476(.A(new_n918_), .B1(G18), .B2(G179), .ZN(new_n919_));
  INV_X1    g0477(.A(new_n919_), .ZN(new_n920_));
  NOR2_X1   g0478(.A1(G18), .A2(G84), .ZN(new_n921_));
  AOI21_X1  g0479(.A(new_n921_), .B1(G18), .B2(G2224), .ZN(new_n922_));
  AOI22_X1  g0480(.A1(new_n915_), .A2(new_n917_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n923_));
  INV_X1    g0481(.A(new_n923_), .ZN(new_n924_));
  OR2_X1    g0482(.A1(new_n920_), .A2(new_n922_), .ZN(new_n925_));
  NOR2_X1   g0483(.A1(G18), .A2(G85), .ZN(new_n926_));
  AOI21_X1  g0484(.A(new_n926_), .B1(G18), .B2(G2230), .ZN(new_n927_));
  INV_X1    g0485(.A(G178), .ZN(new_n928_));
  OAI21_X1  g0486(.A(new_n731_), .B1(new_n507_), .B2(new_n928_), .ZN(new_n929_));
  XOR2_X1   g0487(.A(new_n927_), .B(new_n929_), .Z(new_n930_));
  NAND3_X1  g0488(.A1(new_n924_), .A2(new_n925_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g0489(.A1(new_n507_), .A2(G65), .ZN(new_n932_));
  OAI21_X1  g0490(.A(new_n932_), .B1(new_n507_), .B2(G2211), .ZN(new_n933_));
  XOR2_X1   g0491(.A(new_n933_), .B(KEYINPUT36), .Z(new_n934_));
  INV_X1    g0492(.A(G171), .ZN(new_n935_));
  OAI21_X1  g0493(.A(new_n749_), .B1(new_n507_), .B2(new_n935_), .ZN(new_n936_));
  NAND3_X1  g0494(.A1(new_n930_), .A2(new_n934_), .A3(new_n936_), .ZN(new_n937_));
  XOR2_X1   g0495(.A(new_n937_), .B(KEYINPUT45), .Z(new_n938_));
  OR2_X1    g0496(.A1(new_n915_), .A2(new_n917_), .ZN(new_n939_));
  NAND4_X1  g0497(.A1(new_n911_), .A2(new_n923_), .A3(new_n939_), .A4(new_n925_), .ZN(new_n940_));
  OAI221_X1 g0498(.A(new_n909_), .B1(new_n912_), .B2(new_n931_), .C1(new_n938_), .C2(new_n940_), .ZN(new_n941_));
  OR2_X1    g0499(.A1(new_n941_), .A2(KEYINPUT46), .ZN(new_n942_));
  NAND2_X1  g0500(.A1(new_n941_), .A2(KEYINPUT46), .ZN(new_n943_));
  NAND2_X1  g0501(.A1(new_n927_), .A2(new_n929_), .ZN(new_n944_));
  OAI211_X1 g0502(.A(new_n942_), .B(new_n943_), .C1(new_n910_), .C2(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g0503(.A(new_n901_), .B(new_n903_), .ZN(new_n946_));
  NOR2_X1   g0504(.A1(new_n899_), .A2(new_n946_), .ZN(new_n947_));
  AOI21_X1  g0505(.A(new_n905_), .B1(new_n945_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g0506(.A1(new_n507_), .A2(G112), .ZN(new_n949_));
  OAI21_X1  g0507(.A(new_n949_), .B1(new_n507_), .B2(G1480), .ZN(new_n950_));
  INV_X1    g0508(.A(KEYINPUT34), .ZN(new_n951_));
  XNOR2_X1  g0509(.A(new_n950_), .B(new_n951_), .ZN(new_n952_));
  OR2_X1    g0510(.A1(new_n507_), .A2(G167), .ZN(new_n953_));
  NAND2_X1  g0511(.A1(new_n953_), .A2(new_n695_), .ZN(new_n954_));
  OAI21_X1  g0512(.A(new_n695_), .B1(new_n507_), .B2(G166), .ZN(new_n955_));
  NAND2_X1  g0513(.A1(G18), .A2(G1486), .ZN(new_n956_));
  OAI21_X1  g0514(.A(new_n956_), .B1(G18), .B2(G88), .ZN(new_n957_));
  OAI22_X1  g0515(.A1(new_n952_), .A2(new_n954_), .B1(new_n955_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g0516(.A(new_n958_), .ZN(new_n959_));
  NAND2_X1  g0517(.A1(new_n955_), .A2(new_n957_), .ZN(new_n960_));
  NAND2_X1  g0518(.A1(new_n952_), .A2(new_n954_), .ZN(new_n961_));
  NAND3_X1  g0519(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  OAI21_X1  g0520(.A(new_n695_), .B1(new_n507_), .B2(G168), .ZN(new_n963_));
  NAND2_X1  g0521(.A1(G18), .A2(G106), .ZN(new_n964_));
  OAI21_X1  g0522(.A(new_n964_), .B1(G18), .B2(G87), .ZN(new_n965_));
  XOR2_X1   g0523(.A(new_n963_), .B(new_n965_), .Z(new_n966_));
  OR2_X1    g0524(.A1(new_n507_), .A2(G169), .ZN(new_n967_));
  NAND2_X1  g0525(.A1(new_n967_), .A2(new_n695_), .ZN(new_n968_));
  NAND2_X1  g0526(.A1(G18), .A2(G1469), .ZN(new_n969_));
  OAI21_X1  g0527(.A(new_n969_), .B1(G18), .B2(G111), .ZN(new_n970_));
  NOR2_X1   g0528(.A1(new_n968_), .A2(new_n970_), .ZN(new_n971_));
  INV_X1    g0529(.A(new_n971_), .ZN(new_n972_));
  NAND2_X1  g0530(.A1(new_n968_), .A2(new_n970_), .ZN(new_n973_));
  NAND3_X1  g0531(.A1(new_n966_), .A2(new_n972_), .A3(new_n973_), .ZN(new_n974_));
  NAND2_X1  g0532(.A1(G18), .A2(G1462), .ZN(new_n975_));
  OAI21_X1  g0533(.A(new_n975_), .B1(G18), .B2(G113), .ZN(new_n976_));
  XNOR2_X1  g0534(.A(new_n976_), .B(new_n685_), .ZN(new_n977_));
  NOR3_X1   g0535(.A1(new_n962_), .A2(new_n974_), .A3(new_n977_), .ZN(new_n978_));
  INV_X1    g0536(.A(G4528), .ZN(new_n979_));
  NOR2_X1   g0537(.A1(new_n979_), .A2(G1455), .ZN(new_n980_));
  XOR2_X1   g0538(.A(new_n980_), .B(KEYINPUT35), .Z(new_n981_));
  NOR3_X1   g0539(.A1(new_n981_), .A2(G2204), .A3(new_n979_), .ZN(new_n982_));
  INV_X1    g0540(.A(G2204), .ZN(new_n983_));
  AOI21_X1  g0541(.A(G38), .B1(new_n983_), .B2(G4528), .ZN(new_n984_));
  AOI22_X1  g0542(.A1(new_n982_), .A2(G38), .B1(new_n981_), .B2(new_n984_), .ZN(new_n985_));
  INV_X1    g0543(.A(new_n985_), .ZN(new_n986_));
  NAND2_X1  g0544(.A1(new_n978_), .A2(new_n986_), .ZN(new_n987_));
  NOR2_X1   g0545(.A1(new_n948_), .A2(new_n987_), .ZN(new_n988_));
  XNOR2_X1  g0546(.A(new_n988_), .B(KEYINPUT48), .ZN(new_n989_));
  NAND2_X1  g0547(.A1(new_n507_), .A2(G62), .ZN(new_n990_));
  OAI21_X1  g0548(.A(new_n990_), .B1(new_n507_), .B2(G4437), .ZN(new_n991_));
  XOR2_X1   g0549(.A(new_n991_), .B(KEYINPUT42), .Z(new_n992_));
  AOI21_X1  g0550(.A(new_n532_), .B1(G18), .B2(G189), .ZN(new_n993_));
  OR2_X1    g0551(.A1(new_n992_), .A2(new_n993_), .ZN(new_n994_));
  AOI21_X1  g0552(.A(new_n508_), .B1(G18), .B2(G190), .ZN(new_n995_));
  INV_X1    g0553(.A(new_n995_), .ZN(new_n996_));
  NOR2_X1   g0554(.A1(G18), .A2(G61), .ZN(new_n997_));
  AOI21_X1  g0555(.A(new_n997_), .B1(G18), .B2(G4432), .ZN(new_n998_));
  INV_X1    g0556(.A(new_n525_), .ZN(new_n999_));
  AOI21_X1  g0557(.A(new_n999_), .B1(G18), .B2(G192), .ZN(new_n1000_));
  NOR2_X1   g0558(.A1(G18), .A2(G79), .ZN(new_n1001_));
  AOI21_X1  g0559(.A(new_n1001_), .B1(G18), .B2(G4420), .ZN(new_n1002_));
  INV_X1    g0560(.A(new_n1002_), .ZN(new_n1003_));
  AOI22_X1  g0561(.A1(new_n996_), .A2(new_n998_), .B1(new_n1000_), .B2(new_n1003_), .ZN(new_n1004_));
  INV_X1    g0562(.A(new_n998_), .ZN(new_n1005_));
  NAND2_X1  g0563(.A1(new_n995_), .A2(new_n1005_), .ZN(new_n1006_));
  INV_X1    g0564(.A(new_n1000_), .ZN(new_n1007_));
  NAND2_X1  g0565(.A1(new_n1007_), .A2(new_n1002_), .ZN(new_n1008_));
  AND4_X1   g0566(.A1(new_n994_), .A2(new_n1004_), .A3(new_n1006_), .A4(new_n1008_), .ZN(new_n1009_));
  AOI21_X1  g0567(.A(new_n513_), .B1(G18), .B2(G191), .ZN(new_n1010_));
  XNOR2_X1  g0568(.A(new_n1010_), .B(KEYINPUT43), .ZN(new_n1011_));
  INV_X1    g0569(.A(new_n1011_), .ZN(new_n1012_));
  NOR2_X1   g0570(.A1(G18), .A2(G60), .ZN(new_n1013_));
  AOI21_X1  g0571(.A(new_n1013_), .B1(G18), .B2(G4427), .ZN(new_n1014_));
  NOR2_X1   g0572(.A1(new_n1012_), .A2(new_n1014_), .ZN(new_n1015_));
  INV_X1    g0573(.A(new_n1015_), .ZN(new_n1016_));
  NAND2_X1  g0574(.A1(new_n992_), .A2(new_n993_), .ZN(new_n1017_));
  NAND2_X1  g0575(.A1(new_n1012_), .A2(new_n1014_), .ZN(new_n1018_));
  NAND4_X1  g0576(.A1(new_n1009_), .A2(new_n1016_), .A3(new_n1017_), .A4(new_n1018_), .ZN(new_n1019_));
  XNOR2_X1  g0577(.A(new_n1019_), .B(KEYINPUT44), .ZN(new_n1020_));
  INV_X1    g0578(.A(new_n1020_), .ZN(new_n1021_));
  INV_X1    g0579(.A(G194), .ZN(new_n1022_));
  OAI21_X1  g0580(.A(new_n566_), .B1(new_n507_), .B2(new_n1022_), .ZN(new_n1023_));
  XNOR2_X1  g0581(.A(new_n1023_), .B(KEYINPUT40), .ZN(new_n1024_));
  OR3_X1    g0582(.A1(new_n507_), .A2(KEYINPUT39), .A3(G4410), .ZN(new_n1025_));
  NAND2_X1  g0583(.A1(new_n507_), .A2(G81), .ZN(new_n1026_));
  OAI21_X1  g0584(.A(KEYINPUT39), .B1(new_n507_), .B2(G4410), .ZN(new_n1027_));
  NAND3_X1  g0585(.A1(new_n1025_), .A2(new_n1026_), .A3(new_n1027_), .ZN(new_n1028_));
  NAND2_X1  g0586(.A1(new_n1024_), .A2(new_n1028_), .ZN(new_n1029_));
  NOR2_X1   g0587(.A1(G18), .A2(G59), .ZN(new_n1030_));
  AOI21_X1  g0588(.A(new_n1030_), .B1(G18), .B2(G4405), .ZN(new_n1031_));
  INV_X1    g0589(.A(new_n1031_), .ZN(new_n1032_));
  NOR2_X1   g0590(.A1(new_n546_), .A2(G18), .ZN(new_n1033_));
  AOI21_X1  g0591(.A(new_n1033_), .B1(G18), .B2(G195), .ZN(new_n1034_));
  NOR2_X1   g0592(.A1(new_n1032_), .A2(new_n1034_), .ZN(new_n1035_));
  INV_X1    g0593(.A(new_n1035_), .ZN(new_n1036_));
  NAND2_X1  g0594(.A1(new_n558_), .A2(G18), .ZN(new_n1037_));
  AOI22_X1  g0595(.A1(new_n1037_), .A2(KEYINPUT41), .B1(new_n507_), .B2(G78), .ZN(new_n1038_));
  OAI21_X1  g0596(.A(new_n1038_), .B1(KEYINPUT41), .B2(new_n1037_), .ZN(new_n1039_));
  NAND2_X1  g0597(.A1(G18), .A2(G196), .ZN(new_n1040_));
  OAI21_X1  g0598(.A(new_n1040_), .B1(new_n556_), .B2(G18), .ZN(new_n1041_));
  OR2_X1    g0599(.A1(new_n1039_), .A2(new_n1041_), .ZN(new_n1042_));
  INV_X1    g0600(.A(new_n1034_), .ZN(new_n1043_));
  OAI21_X1  g0601(.A(new_n1042_), .B1(new_n1043_), .B2(new_n1031_), .ZN(new_n1044_));
  INV_X1    g0602(.A(new_n550_), .ZN(new_n1045_));
  AOI21_X1  g0603(.A(new_n1045_), .B1(G18), .B2(G187), .ZN(new_n1046_));
  INV_X1    g0604(.A(new_n1046_), .ZN(new_n1047_));
  NOR2_X1   g0605(.A1(G18), .A2(G77), .ZN(new_n1048_));
  AOI21_X1  g0606(.A(new_n1048_), .B1(G18), .B2(G4394), .ZN(new_n1049_));
  AOI22_X1  g0607(.A1(new_n1047_), .A2(new_n1049_), .B1(new_n1039_), .B2(new_n1041_), .ZN(new_n1050_));
  OAI211_X1 g0608(.A(new_n1029_), .B(new_n1036_), .C1(new_n1044_), .C2(new_n1050_), .ZN(new_n1051_));
  OR2_X1    g0609(.A1(new_n1024_), .A2(new_n1028_), .ZN(new_n1052_));
  NOR2_X1   g0610(.A1(new_n539_), .A2(G18), .ZN(new_n1053_));
  AOI21_X1  g0611(.A(new_n1053_), .B1(G18), .B2(G193), .ZN(new_n1054_));
  INV_X1    g0612(.A(new_n1054_), .ZN(new_n1055_));
  NOR2_X1   g0613(.A1(G18), .A2(G80), .ZN(new_n1056_));
  AOI21_X1  g0614(.A(new_n1056_), .B1(G18), .B2(G4415), .ZN(new_n1057_));
  OR2_X1    g0615(.A1(new_n1055_), .A2(new_n1057_), .ZN(new_n1058_));
  NAND3_X1  g0616(.A1(new_n1051_), .A2(new_n1052_), .A3(new_n1058_), .ZN(new_n1059_));
  NAND2_X1  g0617(.A1(new_n1059_), .A2(KEYINPUT51), .ZN(new_n1060_));
  AND2_X1   g0618(.A1(new_n1052_), .A2(new_n1029_), .ZN(new_n1061_));
  INV_X1    g0619(.A(KEYINPUT51), .ZN(new_n1062_));
  NAND4_X1  g0620(.A1(new_n1061_), .A2(new_n1062_), .A3(new_n1035_), .A4(new_n1058_), .ZN(new_n1063_));
  AOI22_X1  g0621(.A1(new_n1060_), .A2(new_n1063_), .B1(new_n1055_), .B2(new_n1057_), .ZN(new_n1064_));
  NOR2_X1   g0622(.A1(new_n1021_), .A2(new_n1064_), .ZN(new_n1065_));
  OAI221_X1 g0623(.A(new_n1018_), .B1(new_n995_), .B2(new_n1005_), .C1(new_n1015_), .C2(new_n1008_), .ZN(new_n1066_));
  NAND3_X1  g0624(.A1(new_n1066_), .A2(new_n1006_), .A3(new_n1017_), .ZN(new_n1067_));
  NAND2_X1  g0625(.A1(new_n1067_), .A2(new_n994_), .ZN(new_n1068_));
  NOR2_X1   g0626(.A1(new_n1065_), .A2(new_n1068_), .ZN(new_n1069_));
  OR2_X1    g0627(.A1(new_n934_), .A2(new_n936_), .ZN(new_n1070_));
  NAND2_X1  g0628(.A1(new_n934_), .A2(new_n936_), .ZN(new_n1071_));
  NAND3_X1  g0629(.A1(new_n1070_), .A2(new_n1071_), .A3(new_n930_), .ZN(new_n1072_));
  NOR2_X1   g0630(.A1(new_n940_), .A2(new_n1072_), .ZN(new_n1073_));
  NAND2_X1  g0631(.A1(new_n1073_), .A2(new_n947_), .ZN(new_n1074_));
  OR2_X1    g0632(.A1(new_n1074_), .A2(new_n987_), .ZN(new_n1075_));
  NOR2_X1   g0633(.A1(new_n1069_), .A2(new_n1075_), .ZN(new_n1076_));
  XOR2_X1   g0634(.A(new_n1076_), .B(KEYINPUT52), .Z(new_n1077_));
  XNOR2_X1  g0635(.A(new_n1054_), .B(new_n1057_), .ZN(new_n1078_));
  INV_X1    g0636(.A(new_n1049_), .ZN(new_n1079_));
  AOI22_X1  g0637(.A1(new_n1046_), .A2(new_n1079_), .B1(new_n1032_), .B2(new_n1034_), .ZN(new_n1080_));
  AND4_X1   g0638(.A1(new_n1042_), .A2(new_n1078_), .A3(new_n1036_), .A4(new_n1080_), .ZN(new_n1081_));
  AND3_X1   g0639(.A1(new_n1061_), .A2(new_n1050_), .A3(new_n1081_), .ZN(new_n1082_));
  INV_X1    g0640(.A(G203), .ZN(new_n1083_));
  OAI21_X1  g0641(.A(new_n611_), .B1(new_n507_), .B2(new_n1083_), .ZN(new_n1084_));
  XOR2_X1   g0642(.A(new_n1084_), .B(KEYINPUT31), .Z(new_n1085_));
  NOR2_X1   g0643(.A1(G18), .A2(G53), .ZN(new_n1086_));
  AOI21_X1  g0644(.A(new_n1086_), .B1(G18), .B2(G3729), .ZN(new_n1087_));
  NOR2_X1   g0645(.A1(new_n1085_), .A2(new_n1087_), .ZN(new_n1088_));
  NOR2_X1   g0646(.A1(G18), .A2(G56), .ZN(new_n1089_));
  AOI21_X1  g0647(.A(new_n1089_), .B1(G18), .B2(G3749), .ZN(new_n1090_));
  INV_X1    g0648(.A(G200), .ZN(new_n1091_));
  OAI21_X1  g0649(.A(new_n593_), .B1(new_n507_), .B2(new_n1091_), .ZN(new_n1092_));
  NOR2_X1   g0650(.A1(new_n1090_), .A2(new_n1092_), .ZN(new_n1093_));
  AOI21_X1  g0651(.A(new_n605_), .B1(G18), .B2(G202), .ZN(new_n1094_));
  INV_X1    g0652(.A(new_n1094_), .ZN(new_n1095_));
  NOR2_X1   g0653(.A1(G18), .A2(G54), .ZN(new_n1096_));
  AOI21_X1  g0654(.A(new_n1096_), .B1(G18), .B2(G3737), .ZN(new_n1097_));
  AOI21_X1  g0655(.A(new_n1093_), .B1(new_n1095_), .B2(new_n1097_), .ZN(new_n1098_));
  NOR2_X1   g0656(.A1(G18), .A2(G55), .ZN(new_n1099_));
  AOI21_X1  g0657(.A(new_n1099_), .B1(G18), .B2(G3743), .ZN(new_n1100_));
  INV_X1    g0658(.A(G201), .ZN(new_n1101_));
  OAI21_X1  g0659(.A(new_n598_), .B1(new_n507_), .B2(new_n1101_), .ZN(new_n1102_));
  NOR2_X1   g0660(.A1(new_n1100_), .A2(new_n1102_), .ZN(new_n1103_));
  INV_X1    g0661(.A(new_n1097_), .ZN(new_n1104_));
  AOI21_X1  g0662(.A(new_n1103_), .B1(new_n1094_), .B2(new_n1104_), .ZN(new_n1105_));
  AOI22_X1  g0663(.A1(new_n1092_), .A2(new_n1090_), .B1(new_n1100_), .B2(new_n1102_), .ZN(new_n1106_));
  NAND3_X1  g0664(.A1(new_n1098_), .A2(new_n1105_), .A3(new_n1106_), .ZN(new_n1107_));
  INV_X1    g0665(.A(G205), .ZN(new_n1108_));
  OAI21_X1  g0666(.A(new_n626_), .B1(new_n507_), .B2(new_n1108_), .ZN(new_n1109_));
  XOR2_X1   g0667(.A(new_n1109_), .B(KEYINPUT32), .Z(new_n1110_));
  NOR2_X1   g0668(.A1(G18), .A2(G75), .ZN(new_n1111_));
  AOI21_X1  g0669(.A(new_n1111_), .B1(G18), .B2(G3717), .ZN(new_n1112_));
  INV_X1    g0670(.A(new_n1112_), .ZN(new_n1113_));
  NAND2_X1  g0671(.A1(new_n1110_), .A2(new_n1113_), .ZN(new_n1114_));
  NOR2_X1   g0672(.A1(new_n1110_), .A2(new_n1113_), .ZN(new_n1115_));
  NAND2_X1  g0673(.A1(G18), .A2(G3705), .ZN(new_n1116_));
  OAI21_X1  g0674(.A(new_n1116_), .B1(G18), .B2(G74), .ZN(new_n1117_));
  INV_X1    g0675(.A(new_n1117_), .ZN(new_n1118_));
  INV_X1    g0676(.A(G207), .ZN(new_n1119_));
  OAI21_X1  g0677(.A(new_n647_), .B1(new_n507_), .B2(new_n1119_), .ZN(new_n1120_));
  NAND2_X1  g0678(.A1(new_n1118_), .A2(new_n1120_), .ZN(new_n1121_));
  NOR2_X1   g0679(.A1(G18), .A2(G76), .ZN(new_n1122_));
  AOI21_X1  g0680(.A(new_n1122_), .B1(G18), .B2(G3711), .ZN(new_n1123_));
  INV_X1    g0681(.A(G206), .ZN(new_n1124_));
  OAI21_X1  g0682(.A(new_n636_), .B1(new_n507_), .B2(new_n1124_), .ZN(new_n1125_));
  NAND2_X1  g0683(.A1(new_n1123_), .A2(new_n1125_), .ZN(new_n1126_));
  NOR2_X1   g0684(.A1(new_n1118_), .A2(new_n1120_), .ZN(new_n1127_));
  NAND3_X1  g0685(.A1(new_n507_), .A2(G41), .A3(G70), .ZN(new_n1128_));
  OAI211_X1 g0686(.A(new_n1121_), .B(new_n1126_), .C1(new_n1127_), .C2(new_n1128_), .ZN(new_n1129_));
  MUX2_X1   g0687(.A(G103), .B(G204), .S(G18), .Z(new_n1130_));
  NOR2_X1   g0688(.A1(G18), .A2(G73), .ZN(new_n1131_));
  AOI21_X1  g0689(.A(new_n1131_), .B1(G18), .B2(G3723), .ZN(new_n1132_));
  NOR2_X1   g0690(.A1(new_n1130_), .A2(new_n1132_), .ZN(new_n1133_));
  OAI221_X1 g0691(.A(new_n1129_), .B1(KEYINPUT33), .B2(new_n1133_), .C1(new_n1125_), .C2(new_n1123_), .ZN(new_n1134_));
  OR2_X1    g0692(.A1(new_n1134_), .A2(KEYINPUT33), .ZN(new_n1135_));
  AOI21_X1  g0693(.A(new_n1133_), .B1(new_n1120_), .B2(new_n1118_), .ZN(new_n1136_));
  AOI21_X1  g0694(.A(new_n1127_), .B1(new_n1125_), .B2(new_n1123_), .ZN(new_n1137_));
  AND2_X1   g0695(.A1(new_n1130_), .A2(new_n1132_), .ZN(new_n1138_));
  NOR2_X1   g0696(.A1(new_n1123_), .A2(new_n1125_), .ZN(new_n1139_));
  NOR2_X1   g0697(.A1(new_n1138_), .A2(new_n1139_), .ZN(new_n1140_));
  NAND2_X1  g0698(.A1(new_n507_), .A2(G41), .ZN(new_n1141_));
  NOR2_X1   g0699(.A1(G18), .A2(G70), .ZN(new_n1142_));
  NAND2_X1  g0700(.A1(new_n1141_), .A2(new_n1142_), .ZN(new_n1143_));
  AND3_X1   g0701(.A1(new_n1143_), .A2(G89), .A3(new_n1128_), .ZN(new_n1144_));
  NAND4_X1  g0702(.A1(new_n1136_), .A2(new_n1137_), .A3(new_n1140_), .A4(new_n1144_), .ZN(new_n1145_));
  AOI21_X1  g0703(.A(new_n1115_), .B1(new_n1135_), .B2(new_n1145_), .ZN(new_n1146_));
  INV_X1    g0704(.A(new_n1115_), .ZN(new_n1147_));
  AOI21_X1  g0705(.A(new_n1133_), .B1(new_n1134_), .B2(new_n1147_), .ZN(new_n1148_));
  OAI21_X1  g0706(.A(new_n1114_), .B1(new_n1146_), .B2(new_n1148_), .ZN(new_n1149_));
  AOI21_X1  g0707(.A(new_n1138_), .B1(new_n1085_), .B2(new_n1087_), .ZN(new_n1150_));
  AOI211_X1 g0708(.A(new_n1088_), .B(new_n1107_), .C1(new_n1149_), .C2(new_n1150_), .ZN(new_n1151_));
  OAI211_X1 g0709(.A(new_n1095_), .B(new_n1097_), .C1(new_n1100_), .C2(new_n1102_), .ZN(new_n1152_));
  AOI21_X1  g0710(.A(new_n1093_), .B1(new_n1152_), .B2(new_n1106_), .ZN(new_n1153_));
  OAI21_X1  g0711(.A(new_n1082_), .B1(new_n1151_), .B2(new_n1153_), .ZN(new_n1154_));
  OR3_X1    g0712(.A1(new_n1154_), .A2(new_n1075_), .A3(new_n1021_), .ZN(new_n1155_));
  NOR2_X1   g0713(.A1(new_n982_), .A2(new_n817_), .ZN(new_n1156_));
  INV_X1    g0714(.A(new_n974_), .ZN(new_n1157_));
  XOR2_X1   g0715(.A(new_n976_), .B(KEYINPUT49), .Z(new_n1158_));
  AND2_X1   g0716(.A1(new_n1158_), .A2(new_n695_), .ZN(new_n1159_));
  AOI22_X1  g0717(.A1(new_n1157_), .A2(new_n1159_), .B1(new_n966_), .B2(new_n971_), .ZN(new_n1160_));
  NOR2_X1   g0718(.A1(new_n1160_), .A2(new_n962_), .ZN(new_n1161_));
  OR2_X1    g0719(.A1(new_n1161_), .A2(KEYINPUT50), .ZN(new_n1162_));
  NAND2_X1  g0720(.A1(new_n1161_), .A2(KEYINPUT50), .ZN(new_n1163_));
  AOI211_X1 g0721(.A(new_n963_), .B(new_n965_), .C1(new_n952_), .C2(new_n954_), .ZN(new_n1164_));
  OAI21_X1  g0722(.A(new_n960_), .B1(new_n1164_), .B2(new_n958_), .ZN(new_n1165_));
  NAND3_X1  g0723(.A1(new_n1162_), .A2(new_n1163_), .A3(new_n1165_), .ZN(new_n1166_));
  AOI21_X1  g0724(.A(new_n1156_), .B1(new_n1166_), .B2(new_n986_), .ZN(new_n1167_));
  NAND4_X1  g0725(.A1(new_n989_), .A2(new_n1077_), .A3(new_n1155_), .A4(new_n1167_), .ZN(G258));
  NAND4_X1  g0726(.A1(new_n989_), .A2(new_n1077_), .A3(new_n1155_), .A4(new_n1167_), .ZN(G264));
  AOI21_X1  g0727(.A(new_n876_), .B1(new_n858_), .B2(new_n825_), .ZN(new_n1170_));
  INV_X1    g0728(.A(new_n666_), .ZN(new_n1171_));
  NAND3_X1  g0729(.A1(new_n668_), .A2(new_n1171_), .A3(new_n635_), .ZN(new_n1172_));
  INV_X1    g0730(.A(new_n670_), .ZN(new_n1173_));
  NOR2_X1   g0731(.A1(new_n1172_), .A2(new_n1173_), .ZN(new_n1174_));
  NAND2_X1  g0732(.A1(new_n1174_), .A2(KEYINPUT55), .ZN(new_n1175_));
  INV_X1    g0733(.A(new_n681_), .ZN(new_n1176_));
  INV_X1    g0734(.A(new_n547_), .ZN(new_n1177_));
  NOR2_X1   g0735(.A1(new_n1177_), .A2(new_n548_), .ZN(new_n1178_));
  NAND2_X1  g0736(.A1(new_n1177_), .A2(new_n548_), .ZN(new_n1179_));
  AOI21_X1  g0737(.A(new_n1178_), .B1(KEYINPUT54), .B2(new_n1179_), .ZN(new_n1180_));
  OR2_X1    g0738(.A1(new_n1179_), .A2(KEYINPUT54), .ZN(new_n1181_));
  NAND2_X1  g0739(.A1(new_n1180_), .A2(new_n1181_), .ZN(new_n1182_));
  NAND2_X1  g0740(.A1(new_n1182_), .A2(new_n569_), .ZN(new_n1183_));
  NOR3_X1   g0741(.A1(new_n1176_), .A2(new_n1183_), .A3(new_n577_), .ZN(new_n1184_));
  NAND3_X1  g0742(.A1(new_n610_), .A2(new_n676_), .A3(new_n603_), .ZN(new_n1185_));
  INV_X1    g0743(.A(new_n1185_), .ZN(new_n1186_));
  NAND4_X1  g0744(.A1(new_n1175_), .A2(new_n1184_), .A3(G4526), .A4(new_n1186_), .ZN(new_n1187_));
  NOR2_X1   g0745(.A1(new_n1174_), .A2(KEYINPUT55), .ZN(new_n1188_));
  OAI21_X1  g0746(.A(new_n582_), .B1(new_n1187_), .B2(new_n1188_), .ZN(new_n1189_));
  AND2_X1   g0747(.A1(new_n588_), .A2(new_n523_), .ZN(new_n1190_));
  NAND2_X1  g0748(.A1(new_n1189_), .A2(new_n1190_), .ZN(new_n1191_));
  INV_X1    g0749(.A(new_n537_), .ZN(new_n1192_));
  NAND2_X1  g0750(.A1(new_n1191_), .A2(new_n1192_), .ZN(new_n1193_));
  OAI211_X1 g0751(.A(new_n621_), .B(KEYINPUT53), .C1(new_n665_), .C2(new_n1185_), .ZN(new_n1194_));
  NAND2_X1  g0752(.A1(new_n1190_), .A2(new_n1184_), .ZN(new_n1195_));
  OAI21_X1  g0753(.A(new_n621_), .B1(new_n665_), .B2(new_n1185_), .ZN(new_n1196_));
  INV_X1    g0754(.A(KEYINPUT53), .ZN(new_n1197_));
  AOI21_X1  g0755(.A(new_n1195_), .B1(new_n1196_), .B2(new_n1197_), .ZN(new_n1198_));
  AOI21_X1  g0756(.A(new_n1193_), .B1(new_n1194_), .B2(new_n1198_), .ZN(new_n1199_));
  NAND3_X1  g0757(.A1(new_n825_), .A2(new_n717_), .A3(new_n769_), .ZN(new_n1200_));
  OAI21_X1  g0758(.A(new_n1170_), .B1(new_n1199_), .B2(new_n1200_), .ZN(G270));
  INV_X1    g0759(.A(new_n504_), .ZN(new_n1202_));
  INV_X1    g0760(.A(new_n635_), .ZN(new_n1203_));
  NAND2_X1  g0761(.A1(new_n656_), .A2(new_n651_), .ZN(new_n1204_));
  NOR4_X1   g0762(.A1(new_n1203_), .A2(new_n645_), .A3(new_n1204_), .A4(new_n505_), .ZN(new_n1205_));
  AOI21_X1  g0763(.A(new_n1202_), .B1(new_n1205_), .B2(KEYINPUT56), .ZN(new_n1206_));
  OAI21_X1  g0764(.A(new_n1206_), .B1(KEYINPUT56), .B2(new_n1205_), .ZN(new_n1207_));
  NAND3_X1  g0765(.A1(new_n1207_), .A2(new_n662_), .A3(new_n661_), .ZN(new_n1208_));
  XNOR2_X1  g0766(.A(new_n1208_), .B(KEYINPUT58), .ZN(new_n1209_));
  XNOR2_X1  g0767(.A(new_n1209_), .B(KEYINPUT57), .ZN(new_n1210_));
  XNOR2_X1  g0768(.A(new_n1210_), .B(new_n670_), .ZN(G388));
  AND2_X1   g0769(.A1(new_n639_), .A2(new_n642_), .ZN(new_n1212_));
  AND2_X1   g0770(.A1(new_n648_), .A2(new_n650_), .ZN(new_n1213_));
  NAND3_X1  g0771(.A1(new_n1213_), .A2(KEYINPUT15), .A3(new_n649_), .ZN(new_n1214_));
  INV_X1    g0772(.A(KEYINPUT15), .ZN(new_n1215_));
  NAND2_X1  g0773(.A1(new_n651_), .A2(new_n1215_), .ZN(new_n1216_));
  AOI21_X1  g0774(.A(new_n1212_), .B1(new_n1214_), .B2(new_n1216_), .ZN(new_n1217_));
  XOR2_X1   g0775(.A(new_n659_), .B(KEYINPUT59), .Z(new_n1218_));
  NOR2_X1   g0776(.A1(new_n1217_), .A2(new_n1218_), .ZN(new_n1219_));
  INV_X1    g0777(.A(new_n1204_), .ZN(new_n1220_));
  NAND2_X1  g0778(.A1(new_n668_), .A2(new_n1220_), .ZN(new_n1221_));
  INV_X1    g0779(.A(new_n503_), .ZN(new_n1222_));
  AOI21_X1  g0780(.A(new_n501_), .B1(new_n1222_), .B2(G4526), .ZN(new_n1223_));
  OAI21_X1  g0781(.A(new_n1219_), .B1(new_n1221_), .B2(new_n1223_), .ZN(new_n1224_));
  XNOR2_X1  g0782(.A(new_n635_), .B(KEYINPUT60), .ZN(new_n1225_));
  XNOR2_X1  g0783(.A(new_n1224_), .B(new_n1225_), .ZN(G391));
  INV_X1    g0784(.A(KEYINPUT61), .ZN(new_n1227_));
  AOI21_X1  g0785(.A(new_n667_), .B1(new_n1227_), .B2(new_n652_), .ZN(new_n1228_));
  INV_X1    g0786(.A(KEYINPUT62), .ZN(new_n1229_));
  AOI21_X1  g0787(.A(new_n654_), .B1(new_n1213_), .B2(new_n1229_), .ZN(new_n1230_));
  OAI21_X1  g0788(.A(new_n1230_), .B1(new_n1229_), .B2(new_n1213_), .ZN(new_n1231_));
  NAND3_X1  g0789(.A1(new_n654_), .A2(new_n655_), .A3(KEYINPUT62), .ZN(new_n1232_));
  NAND3_X1  g0790(.A1(new_n1231_), .A2(new_n501_), .A3(new_n1232_), .ZN(new_n1233_));
  OAI211_X1 g0791(.A(new_n1228_), .B(new_n1233_), .C1(new_n1227_), .C2(new_n652_), .ZN(new_n1234_));
  XNOR2_X1  g0792(.A(new_n1212_), .B(KEYINPUT63), .ZN(new_n1235_));
  XNOR2_X1  g0793(.A(new_n1234_), .B(new_n1235_), .ZN(G394));
  XOR2_X1   g0794(.A(new_n1204_), .B(new_n1223_), .Z(G397));
  NAND2_X1  g0795(.A1(new_n609_), .A2(new_n674_), .ZN(new_n1238_));
  NAND2_X1  g0796(.A1(new_n1238_), .A2(new_n608_), .ZN(new_n1239_));
  AND2_X1   g0797(.A1(new_n1239_), .A2(new_n603_), .ZN(new_n1240_));
  OR2_X1    g0798(.A1(new_n1240_), .A2(new_n617_), .ZN(new_n1241_));
  NAND2_X1  g0799(.A1(new_n672_), .A2(new_n1241_), .ZN(new_n1242_));
  INV_X1    g0800(.A(KEYINPUT64), .ZN(new_n1243_));
  AND2_X1   g0801(.A1(new_n616_), .A2(new_n1243_), .ZN(new_n1244_));
  NOR2_X1   g0802(.A1(new_n616_), .A2(new_n1243_), .ZN(new_n1245_));
  OAI21_X1  g0803(.A(new_n618_), .B1(new_n1244_), .B2(new_n1245_), .ZN(new_n1246_));
  XNOR2_X1  g0804(.A(new_n1246_), .B(KEYINPUT65), .ZN(new_n1247_));
  OAI21_X1  g0805(.A(new_n1242_), .B1(new_n1247_), .B2(new_n672_), .ZN(new_n1248_));
  XNOR2_X1  g0806(.A(new_n1248_), .B(new_n673_), .ZN(G376));
  NAND2_X1  g0807(.A1(new_n615_), .A2(new_n609_), .ZN(new_n1250_));
  NAND2_X1  g0808(.A1(new_n1250_), .A2(new_n608_), .ZN(new_n1251_));
  XOR2_X1   g0809(.A(new_n604_), .B(new_n1251_), .Z(new_n1252_));
  NOR2_X1   g0810(.A1(new_n672_), .A2(new_n1252_), .ZN(new_n1253_));
  XNOR2_X1  g0811(.A(new_n1239_), .B(new_n603_), .ZN(new_n1254_));
  AOI21_X1  g0812(.A(new_n1253_), .B1(new_n672_), .B2(new_n1254_), .ZN(G379));
  AOI21_X1  g0813(.A(new_n615_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n1256_));
  XNOR2_X1  g0814(.A(new_n1256_), .B(new_n610_), .ZN(G382));
  XNOR2_X1  g0815(.A(new_n675_), .B(KEYINPUT66), .ZN(new_n1258_));
  XNOR2_X1  g0816(.A(new_n672_), .B(new_n1258_), .ZN(G385));
  NAND2_X1  g0817(.A1(new_n749_), .A2(new_n742_), .ZN(new_n1260_));
  NAND2_X1  g0818(.A1(new_n719_), .A2(new_n720_), .ZN(new_n1261_));
  XNOR2_X1  g0819(.A(new_n1260_), .B(new_n1261_), .ZN(new_n1262_));
  NAND2_X1  g0820(.A1(new_n507_), .A2(G141), .ZN(new_n1263_));
  INV_X1    g0821(.A(new_n1263_), .ZN(new_n1264_));
  AOI21_X1  g0822(.A(new_n1264_), .B1(G18), .B2(G161), .ZN(new_n1265_));
  XNOR2_X1  g0823(.A(new_n1262_), .B(new_n1265_), .ZN(new_n1266_));
  XNOR2_X1  g0824(.A(new_n1266_), .B(new_n853_), .ZN(new_n1267_));
  XNOR2_X1  g0825(.A(new_n761_), .B(new_n753_), .ZN(new_n1268_));
  XNOR2_X1  g0826(.A(new_n1268_), .B(new_n687_), .ZN(new_n1269_));
  XNOR2_X1  g0827(.A(new_n1267_), .B(new_n1269_), .ZN(new_n1270_));
  OR2_X1    g0828(.A1(new_n507_), .A2(G155), .ZN(new_n1271_));
  OAI22_X1  g0829(.A1(new_n700_), .A2(new_n1271_), .B1(new_n694_), .B2(new_n711_), .ZN(new_n1272_));
  XOR2_X1   g0830(.A(new_n1272_), .B(new_n706_), .Z(new_n1273_));
  NOR2_X1   g0831(.A1(new_n1270_), .A2(new_n1273_), .ZN(new_n1274_));
  NAND2_X1  g0832(.A1(new_n1270_), .A2(new_n1273_), .ZN(new_n1275_));
  INV_X1    g0833(.A(G229), .ZN(new_n1276_));
  OAI21_X1  g0834(.A(new_n1141_), .B1(new_n507_), .B2(new_n1276_), .ZN(new_n1277_));
  XNOR2_X1  g0835(.A(new_n1213_), .B(new_n1277_), .ZN(new_n1278_));
  XNOR2_X1  g0836(.A(new_n1278_), .B(new_n613_), .ZN(new_n1279_));
  XNOR2_X1  g0837(.A(new_n606_), .B(new_n595_), .ZN(new_n1280_));
  XNOR2_X1  g0838(.A(new_n1280_), .B(new_n600_), .ZN(new_n1281_));
  XNOR2_X1  g0839(.A(new_n1279_), .B(new_n1281_), .ZN(new_n1282_));
  XOR2_X1   g0840(.A(new_n628_), .B(new_n638_), .Z(new_n1283_));
  XNOR2_X1  g0841(.A(new_n1283_), .B(new_n624_), .ZN(new_n1284_));
  NAND2_X1  g0842(.A1(new_n507_), .A2(G44), .ZN(new_n1285_));
  INV_X1    g0843(.A(G239), .ZN(new_n1286_));
  OAI21_X1  g0844(.A(new_n1285_), .B1(new_n507_), .B2(new_n1286_), .ZN(new_n1287_));
  XOR2_X1   g0845(.A(new_n1284_), .B(new_n1287_), .Z(new_n1288_));
  XNOR2_X1  g0846(.A(new_n1282_), .B(new_n1288_), .ZN(new_n1289_));
  OAI21_X1  g0847(.A(new_n791_), .B1(new_n507_), .B2(G215), .ZN(new_n1290_));
  OAI21_X1  g0848(.A(new_n1290_), .B1(new_n781_), .B2(new_n791_), .ZN(new_n1291_));
  NAND3_X1  g0849(.A1(new_n773_), .A2(G18), .A3(new_n805_), .ZN(new_n1292_));
  NAND3_X1  g0850(.A1(new_n806_), .A2(G18), .A3(new_n772_), .ZN(new_n1293_));
  NAND2_X1  g0851(.A1(new_n1292_), .A2(new_n1293_), .ZN(new_n1294_));
  XNOR2_X1  g0852(.A(new_n1291_), .B(new_n1294_), .ZN(new_n1295_));
  NOR2_X1   g0853(.A1(new_n1295_), .A2(KEYINPUT67), .ZN(new_n1296_));
  NOR3_X1   g0854(.A1(new_n685_), .A2(new_n507_), .A3(G209), .ZN(new_n1297_));
  XNOR2_X1  g0855(.A(new_n1296_), .B(new_n1297_), .ZN(new_n1298_));
  NAND2_X1  g0856(.A1(new_n695_), .A2(G18), .ZN(new_n1299_));
  INV_X1    g0857(.A(G211), .ZN(new_n1300_));
  OR2_X1    g0858(.A1(new_n1300_), .A2(G212), .ZN(new_n1301_));
  NAND2_X1  g0859(.A1(new_n1300_), .A2(G212), .ZN(new_n1302_));
  AOI21_X1  g0860(.A(new_n1299_), .B1(new_n1301_), .B2(new_n1302_), .ZN(new_n1303_));
  XNOR2_X1  g0861(.A(new_n1298_), .B(new_n1303_), .ZN(new_n1304_));
  NAND3_X1  g0862(.A1(new_n1275_), .A2(new_n1289_), .A3(new_n1304_), .ZN(new_n1305_));
  XNOR2_X1  g0863(.A(new_n547_), .B(new_n557_), .ZN(new_n1306_));
  XOR2_X1   g0864(.A(new_n1306_), .B(KEYINPUT69), .Z(new_n1307_));
  INV_X1    g0865(.A(new_n1307_), .ZN(new_n1308_));
  XNOR2_X1  g0866(.A(new_n568_), .B(new_n540_), .ZN(new_n1309_));
  XOR2_X1   g0867(.A(new_n1309_), .B(KEYINPUT68), .Z(new_n1310_));
  NAND2_X1  g0868(.A1(new_n507_), .A2(G115), .ZN(new_n1311_));
  INV_X1    g0869(.A(G227), .ZN(new_n1312_));
  OAI21_X1  g0870(.A(new_n1311_), .B1(new_n507_), .B2(new_n1312_), .ZN(new_n1313_));
  XNOR2_X1  g0871(.A(new_n552_), .B(new_n1313_), .ZN(new_n1314_));
  INV_X1    g0872(.A(new_n1314_), .ZN(new_n1315_));
  NAND3_X1  g0873(.A1(new_n1308_), .A2(new_n1310_), .A3(new_n1315_), .ZN(new_n1316_));
  XNOR2_X1  g0874(.A(new_n1316_), .B(KEYINPUT70), .ZN(new_n1317_));
  NAND2_X1  g0875(.A1(new_n1307_), .A2(new_n1314_), .ZN(new_n1318_));
  NAND3_X1  g0876(.A1(new_n1318_), .A2(new_n1309_), .A3(new_n1306_), .ZN(new_n1319_));
  AOI22_X1  g0877(.A1(new_n1318_), .A2(new_n1309_), .B1(new_n1310_), .B2(new_n1306_), .ZN(new_n1320_));
  OAI211_X1 g0878(.A(new_n1317_), .B(new_n1319_), .C1(new_n1315_), .C2(new_n1320_), .ZN(new_n1321_));
  INV_X1    g0879(.A(new_n527_), .ZN(new_n1322_));
  XNOR2_X1  g0880(.A(new_n1322_), .B(new_n533_), .ZN(new_n1323_));
  XNOR2_X1  g0881(.A(new_n1323_), .B(new_n509_), .ZN(new_n1324_));
  XNOR2_X1  g0882(.A(new_n1321_), .B(new_n1324_), .ZN(new_n1325_));
  XNOR2_X1  g0883(.A(new_n521_), .B(KEYINPUT71), .ZN(new_n1326_));
  AOI211_X1 g0884(.A(new_n1274_), .B(new_n1305_), .C1(new_n1325_), .C2(new_n1326_), .ZN(new_n1327_));
  OAI21_X1  g0885(.A(new_n1327_), .B1(new_n1326_), .B2(new_n1325_), .ZN(G412));
  XNOR2_X1  g0886(.A(new_n1118_), .B(new_n1132_), .ZN(new_n1329_));
  XNOR2_X1  g0887(.A(new_n1329_), .B(new_n1123_), .ZN(new_n1330_));
  NAND2_X1  g0888(.A1(new_n507_), .A2(G69), .ZN(new_n1331_));
  OAI21_X1  g0889(.A(new_n1331_), .B1(new_n507_), .B2(G3698), .ZN(new_n1332_));
  XNOR2_X1  g0890(.A(new_n1330_), .B(new_n1332_), .ZN(new_n1333_));
  AOI21_X1  g0891(.A(new_n1142_), .B1(G18), .B2(G3701), .ZN(new_n1334_));
  XNOR2_X1  g0892(.A(new_n1112_), .B(new_n1334_), .ZN(new_n1335_));
  XNOR2_X1  g0893(.A(new_n1333_), .B(new_n1335_), .ZN(new_n1336_));
  XNOR2_X1  g0894(.A(new_n1100_), .B(new_n1097_), .ZN(new_n1337_));
  XNOR2_X1  g0895(.A(new_n1336_), .B(new_n1337_), .ZN(new_n1338_));
  XNOR2_X1  g0896(.A(new_n1090_), .B(new_n1087_), .ZN(new_n1339_));
  XNOR2_X1  g0897(.A(new_n1338_), .B(new_n1339_), .ZN(new_n1340_));
  NAND2_X1  g0898(.A1(G18), .A2(G2208), .ZN(new_n1341_));
  OAI21_X1  g0899(.A(new_n1341_), .B1(G18), .B2(G82), .ZN(new_n1342_));
  XNOR2_X1  g0900(.A(new_n922_), .B(new_n1342_), .ZN(new_n1343_));
  XNOR2_X1  g0901(.A(new_n1343_), .B(new_n917_), .ZN(new_n1344_));
  OR2_X1    g0902(.A1(new_n1344_), .A2(new_n934_), .ZN(new_n1345_));
  NAND2_X1  g0903(.A1(new_n1344_), .A2(new_n934_), .ZN(new_n1346_));
  NAND3_X1  g0904(.A1(new_n1345_), .A2(KEYINPUT72), .A3(new_n1346_), .ZN(new_n1347_));
  XNOR2_X1  g0905(.A(new_n881_), .B(new_n903_), .ZN(new_n1348_));
  XNOR2_X1  g0906(.A(new_n927_), .B(new_n908_), .ZN(new_n1349_));
  XNOR2_X1  g0907(.A(new_n1348_), .B(new_n1349_), .ZN(new_n1350_));
  XNOR2_X1  g0908(.A(new_n1347_), .B(new_n1350_), .ZN(new_n1351_));
  XOR2_X1   g0909(.A(new_n888_), .B(new_n891_), .Z(new_n1352_));
  XNOR2_X1  g0910(.A(new_n1351_), .B(new_n1352_), .ZN(new_n1353_));
  XOR2_X1   g0911(.A(new_n1002_), .B(new_n1014_), .Z(new_n1354_));
  XNOR2_X1  g0912(.A(new_n1354_), .B(new_n992_), .ZN(new_n1355_));
  NAND2_X1  g0913(.A1(G18), .A2(G4393), .ZN(new_n1356_));
  OAI21_X1  g0914(.A(new_n1356_), .B1(G18), .B2(G58), .ZN(new_n1357_));
  XNOR2_X1  g0915(.A(new_n1057_), .B(new_n1357_), .ZN(new_n1358_));
  XNOR2_X1  g0916(.A(new_n1358_), .B(new_n1005_), .ZN(new_n1359_));
  XNOR2_X1  g0917(.A(new_n1355_), .B(new_n1359_), .ZN(new_n1360_));
  XOR2_X1   g0918(.A(new_n1049_), .B(new_n1031_), .Z(new_n1361_));
  XNOR2_X1  g0919(.A(new_n1361_), .B(new_n1039_), .ZN(new_n1362_));
  XNOR2_X1  g0920(.A(new_n1362_), .B(new_n1028_), .ZN(new_n1363_));
  XNOR2_X1  g0921(.A(new_n1360_), .B(new_n1363_), .ZN(new_n1364_));
  XOR2_X1   g0922(.A(new_n952_), .B(new_n957_), .Z(new_n1365_));
  XOR2_X1   g0923(.A(new_n965_), .B(new_n970_), .Z(new_n1366_));
  OR2_X1    g0924(.A1(new_n1365_), .A2(new_n1366_), .ZN(new_n1367_));
  NAND2_X1  g0925(.A1(new_n1365_), .A2(new_n1366_), .ZN(new_n1368_));
  NAND2_X1  g0926(.A1(new_n507_), .A2(G114), .ZN(new_n1369_));
  OAI21_X1  g0927(.A(new_n1369_), .B1(new_n507_), .B2(G1459), .ZN(new_n1370_));
  XNOR2_X1  g0928(.A(new_n1158_), .B(new_n1370_), .ZN(new_n1371_));
  NAND3_X1  g0929(.A1(new_n1367_), .A2(new_n1368_), .A3(new_n1371_), .ZN(new_n1372_));
  NOR2_X1   g0930(.A1(new_n1368_), .A2(new_n1371_), .ZN(new_n1373_));
  AND2_X1   g0931(.A1(new_n1373_), .A2(KEYINPUT73), .ZN(new_n1374_));
  NOR2_X1   g0932(.A1(new_n1373_), .A2(KEYINPUT73), .ZN(new_n1375_));
  OAI221_X1 g0933(.A(new_n1372_), .B1(new_n1371_), .B2(new_n1367_), .C1(new_n1374_), .C2(new_n1375_), .ZN(new_n1376_));
  NAND2_X1  g0934(.A1(new_n507_), .A2(G1455), .ZN(new_n1377_));
  OAI21_X1  g0935(.A(new_n1377_), .B1(new_n507_), .B2(G1492), .ZN(new_n1378_));
  XNOR2_X1  g0936(.A(new_n1376_), .B(new_n1378_), .ZN(new_n1379_));
  NAND2_X1  g0937(.A1(G18), .A2(G1496), .ZN(new_n1380_));
  OAI21_X1  g0938(.A(new_n1380_), .B1(G18), .B2(G2204), .ZN(new_n1381_));
  OAI211_X1 g0939(.A(new_n1353_), .B(new_n1364_), .C1(new_n1379_), .C2(new_n1381_), .ZN(new_n1382_));
  AOI211_X1 g0940(.A(new_n1340_), .B(new_n1382_), .C1(new_n1381_), .C2(new_n1379_), .ZN(new_n1383_));
  XOR2_X1   g0941(.A(new_n1383_), .B(KEYINPUT74), .Z(G414));
  XNOR2_X1  g0942(.A(new_n1024_), .B(new_n1047_), .ZN(new_n1385_));
  INV_X1    g0943(.A(new_n1311_), .ZN(new_n1386_));
  AOI21_X1  g0944(.A(new_n1386_), .B1(G18), .B2(G197), .ZN(new_n1387_));
  XNOR2_X1  g0945(.A(new_n1385_), .B(new_n1387_), .ZN(new_n1388_));
  XNOR2_X1  g0946(.A(new_n1388_), .B(new_n1043_), .ZN(new_n1389_));
  XOR2_X1   g0947(.A(new_n1054_), .B(KEYINPUT78), .Z(new_n1390_));
  XNOR2_X1  g0948(.A(new_n1390_), .B(new_n1041_), .ZN(new_n1391_));
  XNOR2_X1  g0949(.A(new_n1391_), .B(new_n1012_), .ZN(new_n1392_));
  XNOR2_X1  g0950(.A(new_n1389_), .B(new_n1392_), .ZN(new_n1393_));
  XOR2_X1   g0951(.A(new_n993_), .B(KEYINPUT79), .Z(new_n1394_));
  XNOR2_X1  g0952(.A(new_n1000_), .B(new_n995_), .ZN(new_n1395_));
  XNOR2_X1  g0953(.A(new_n1394_), .B(new_n1395_), .ZN(new_n1396_));
  AND2_X1   g0954(.A1(new_n1393_), .A2(new_n1396_), .ZN(new_n1397_));
  NOR2_X1   g0955(.A1(new_n1393_), .A2(new_n1396_), .ZN(new_n1398_));
  MUX2_X1   g0956(.A(new_n953_), .B(new_n954_), .S(new_n955_), .Z(new_n1399_));
  MUX2_X1   g0957(.A(new_n967_), .B(new_n968_), .S(new_n963_), .Z(new_n1400_));
  XNOR2_X1  g0958(.A(new_n1399_), .B(new_n1400_), .ZN(new_n1401_));
  NOR2_X1   g0959(.A1(new_n1299_), .A2(G170), .ZN(new_n1402_));
  XNOR2_X1  g0960(.A(new_n1402_), .B(KEYINPUT80), .ZN(new_n1403_));
  XNOR2_X1  g0961(.A(G164), .B(G165), .ZN(new_n1404_));
  NOR2_X1   g0962(.A1(new_n1404_), .A2(new_n1299_), .ZN(new_n1405_));
  XNOR2_X1  g0963(.A(new_n1403_), .B(new_n1405_), .ZN(new_n1406_));
  XNOR2_X1  g0964(.A(new_n1401_), .B(new_n1406_), .ZN(new_n1407_));
  NOR3_X1   g0965(.A1(new_n1397_), .A2(new_n1398_), .A3(new_n1407_), .ZN(new_n1408_));
  INV_X1    g0966(.A(G198), .ZN(new_n1409_));
  OAI21_X1  g0967(.A(new_n1141_), .B1(new_n507_), .B2(new_n1409_), .ZN(new_n1410_));
  INV_X1    g0968(.A(G208), .ZN(new_n1411_));
  OAI21_X1  g0969(.A(new_n1285_), .B1(new_n507_), .B2(new_n1411_), .ZN(new_n1412_));
  XOR2_X1   g0970(.A(new_n1410_), .B(new_n1412_), .Z(new_n1413_));
  XNOR2_X1  g0971(.A(new_n1130_), .B(new_n1109_), .ZN(new_n1414_));
  OR2_X1    g0972(.A1(new_n1413_), .A2(new_n1414_), .ZN(new_n1415_));
  XOR2_X1   g0973(.A(new_n1120_), .B(new_n1125_), .Z(new_n1416_));
  NOR2_X1   g0974(.A1(new_n1415_), .A2(new_n1416_), .ZN(new_n1417_));
  XOR2_X1   g0975(.A(new_n1417_), .B(KEYINPUT76), .Z(new_n1418_));
  NAND2_X1  g0976(.A1(new_n1413_), .A2(new_n1414_), .ZN(new_n1419_));
  NOR2_X1   g0977(.A1(new_n1419_), .A2(new_n1416_), .ZN(new_n1420_));
  XOR2_X1   g0978(.A(new_n1420_), .B(KEYINPUT75), .Z(new_n1421_));
  NAND3_X1  g0979(.A1(new_n1415_), .A2(new_n1416_), .A3(new_n1419_), .ZN(new_n1422_));
  NAND3_X1  g0980(.A1(new_n1418_), .A2(new_n1421_), .A3(new_n1422_), .ZN(new_n1423_));
  XNOR2_X1  g0981(.A(new_n1094_), .B(new_n1102_), .ZN(new_n1424_));
  XOR2_X1   g0982(.A(new_n1424_), .B(new_n1085_), .Z(new_n1425_));
  XNOR2_X1  g0983(.A(new_n1423_), .B(new_n1425_), .ZN(new_n1426_));
  XOR2_X1   g0984(.A(new_n1092_), .B(KEYINPUT77), .Z(new_n1427_));
  XNOR2_X1  g0985(.A(new_n1426_), .B(new_n1427_), .ZN(new_n1428_));
  XNOR2_X1  g0986(.A(new_n936_), .B(new_n929_), .ZN(new_n1429_));
  XNOR2_X1  g0987(.A(new_n1429_), .B(new_n906_), .ZN(new_n1430_));
  XNOR2_X1  g0988(.A(new_n1430_), .B(new_n920_), .ZN(new_n1431_));
  MUX2_X1   g0989(.A(new_n885_), .B(new_n886_), .S(new_n900_), .Z(new_n1432_));
  XNOR2_X1  g0990(.A(new_n1432_), .B(new_n879_), .ZN(new_n1433_));
  XNOR2_X1  g0991(.A(new_n1431_), .B(new_n1433_), .ZN(new_n1434_));
  AOI21_X1  g0992(.A(new_n1264_), .B1(G18), .B2(G181), .ZN(new_n1435_));
  XOR2_X1   g0993(.A(new_n914_), .B(new_n1435_), .Z(new_n1436_));
  XNOR2_X1  g0994(.A(new_n1436_), .B(new_n893_), .ZN(new_n1437_));
  XNOR2_X1  g0995(.A(new_n1434_), .B(new_n1437_), .ZN(new_n1438_));
  NAND3_X1  g0996(.A1(new_n1408_), .A2(new_n1428_), .A3(new_n1438_), .ZN(G416));
  NAND2_X1  g0997(.A1(new_n1154_), .A2(new_n1064_), .ZN(new_n1440_));
  AOI21_X1  g0998(.A(new_n1068_), .B1(new_n1440_), .B2(new_n1020_), .ZN(new_n1441_));
  OAI21_X1  g0999(.A(new_n948_), .B1(new_n1441_), .B2(new_n1074_), .ZN(new_n1442_));
  AOI21_X1  g1000(.A(new_n1166_), .B1(new_n1442_), .B2(new_n978_), .ZN(new_n1443_));
  OAI22_X1  g1001(.A1(new_n1443_), .A2(new_n985_), .B1(new_n817_), .B2(new_n982_), .ZN(new_n1444_));
  XNOR2_X1  g1002(.A(new_n1444_), .B(KEYINPUT81), .ZN(G249));
  NOR2_X1   g1003(.A1(new_n748_), .A2(new_n750_), .ZN(new_n1446_));
  XNOR2_X1  g1004(.A(new_n684_), .B(new_n1446_), .ZN(G295));
  NOR2_X1   g1005(.A1(new_n771_), .A2(new_n858_), .ZN(new_n1448_));
  XNOR2_X1  g1006(.A(new_n1448_), .B(new_n803_), .ZN(new_n1449_));
  XNOR2_X1  g1007(.A(new_n1449_), .B(KEYINPUT82), .ZN(G324));
  XNOR2_X1  g1008(.A(new_n1441_), .B(KEYINPUT83), .ZN(G252));
  AND3_X1   g1009(.A1(new_n1196_), .A2(new_n1190_), .A3(new_n1184_), .ZN(new_n1452_));
  OAI211_X1 g1010(.A(new_n717_), .B(new_n769_), .C1(new_n1452_), .C2(new_n1193_), .ZN(new_n1453_));
  XNOR2_X1  g1011(.A(new_n858_), .B(KEYINPUT84), .ZN(new_n1454_));
  NAND2_X1  g1012(.A1(new_n1453_), .A2(new_n1454_), .ZN(new_n1455_));
  AOI21_X1  g1013(.A(new_n874_), .B1(new_n1455_), .B2(new_n813_), .ZN(new_n1456_));
  OAI21_X1  g1014(.A(new_n862_), .B1(new_n1456_), .B2(new_n824_), .ZN(G276));
  NOR2_X1   g1015(.A1(new_n848_), .A2(new_n722_), .ZN(new_n1458_));
  INV_X1    g1016(.A(new_n1458_), .ZN(new_n1459_));
  AOI21_X1  g1017(.A(new_n854_), .B1(new_n740_), .B2(new_n835_), .ZN(new_n1460_));
  NAND2_X1  g1018(.A1(new_n734_), .A2(new_n739_), .ZN(new_n1461_));
  NAND4_X1  g1019(.A1(new_n1461_), .A2(new_n839_), .A3(new_n750_), .A4(new_n841_), .ZN(new_n1462_));
  NAND3_X1  g1020(.A1(new_n1459_), .A2(new_n1460_), .A3(new_n1462_), .ZN(new_n1463_));
  INV_X1    g1021(.A(new_n1463_), .ZN(new_n1464_));
  INV_X1    g1022(.A(new_n1446_), .ZN(new_n1465_));
  NOR2_X1   g1023(.A1(new_n684_), .A2(new_n1465_), .ZN(new_n1466_));
  NAND3_X1  g1024(.A1(new_n1466_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n1467_));
  OAI21_X1  g1025(.A(new_n1464_), .B1(new_n1467_), .B2(new_n848_), .ZN(new_n1468_));
  XNOR2_X1  g1026(.A(new_n1468_), .B(new_n768_), .ZN(G310));
  OAI211_X1 g1027(.A(new_n836_), .B(new_n842_), .C1(new_n1467_), .C2(KEYINPUT85), .ZN(new_n1470_));
  AOI21_X1  g1028(.A(new_n1470_), .B1(KEYINPUT85), .B2(new_n1467_), .ZN(new_n1471_));
  XNOR2_X1  g1029(.A(new_n1471_), .B(new_n1461_), .ZN(G313));
  NAND2_X1  g1030(.A1(new_n755_), .A2(KEYINPUT20), .ZN(new_n1473_));
  INV_X1    g1031(.A(KEYINPUT86), .ZN(new_n1474_));
  NAND2_X1  g1032(.A1(new_n838_), .A2(new_n833_), .ZN(new_n1475_));
  NAND3_X1  g1033(.A1(new_n1473_), .A2(new_n1474_), .A3(new_n1475_), .ZN(new_n1476_));
  OAI21_X1  g1034(.A(KEYINPUT86), .B1(new_n832_), .B2(new_n834_), .ZN(new_n1477_));
  NAND2_X1  g1035(.A1(new_n1260_), .A2(new_n741_), .ZN(new_n1478_));
  OAI211_X1 g1036(.A(new_n1476_), .B(new_n1477_), .C1(new_n758_), .C2(new_n1478_), .ZN(new_n1479_));
  AOI21_X1  g1037(.A(new_n1479_), .B1(new_n1466_), .B2(new_n839_), .ZN(new_n1480_));
  XNOR2_X1  g1038(.A(new_n1480_), .B(new_n841_), .ZN(G316));
  NOR2_X1   g1039(.A1(new_n1466_), .A2(new_n750_), .ZN(new_n1482_));
  XNOR2_X1  g1040(.A(new_n1482_), .B(new_n839_), .ZN(G319));
  NOR2_X1   g1041(.A1(new_n1448_), .A2(new_n804_), .ZN(new_n1484_));
  XNOR2_X1  g1042(.A(new_n800_), .B(KEYINPUT87), .ZN(new_n1485_));
  NAND2_X1  g1043(.A1(new_n1485_), .A2(new_n796_), .ZN(new_n1486_));
  NAND2_X1  g1044(.A1(new_n1486_), .A2(new_n867_), .ZN(new_n1487_));
  AOI21_X1  g1045(.A(new_n872_), .B1(new_n1487_), .B2(new_n789_), .ZN(new_n1488_));
  INV_X1    g1046(.A(new_n1488_), .ZN(new_n1489_));
  NOR2_X1   g1047(.A1(new_n1484_), .A2(new_n1489_), .ZN(new_n1490_));
  XNOR2_X1  g1048(.A(new_n1490_), .B(new_n811_), .ZN(G327));
  NAND2_X1  g1049(.A1(new_n868_), .A2(new_n787_), .ZN(new_n1492_));
  OAI21_X1  g1050(.A(new_n803_), .B1(new_n771_), .B2(new_n858_), .ZN(new_n1493_));
  NAND2_X1  g1051(.A1(new_n796_), .A2(new_n787_), .ZN(new_n1494_));
  OAI211_X1 g1052(.A(new_n871_), .B(new_n1492_), .C1(new_n1493_), .C2(new_n1494_), .ZN(new_n1495_));
  XNOR2_X1  g1053(.A(new_n1495_), .B(new_n779_), .ZN(G330));
  INV_X1    g1054(.A(new_n1485_), .ZN(new_n1497_));
  AND2_X1   g1055(.A1(new_n1493_), .A2(new_n1497_), .ZN(new_n1498_));
  OAI21_X1  g1056(.A(new_n793_), .B1(new_n1498_), .B2(new_n795_), .ZN(new_n1499_));
  NAND2_X1  g1057(.A1(new_n1499_), .A2(new_n788_), .ZN(new_n1500_));
  OAI211_X1 g1058(.A(new_n787_), .B(new_n793_), .C1(new_n1498_), .C2(new_n795_), .ZN(new_n1501_));
  NAND2_X1  g1059(.A1(new_n1500_), .A2(new_n1501_), .ZN(G333));
  XNOR2_X1  g1060(.A(new_n1498_), .B(new_n796_), .ZN(G336));
  NOR4_X1   g1061(.A1(G404), .A2(G406), .A3(G408), .A4(G410), .ZN(new_n1504_));
  XNOR2_X1  g1062(.A(new_n1383_), .B(KEYINPUT74), .ZN(new_n1505_));
  INV_X1    g1063(.A(KEYINPUT88), .ZN(new_n1506_));
  NOR2_X1   g1064(.A1(G412), .A2(G416), .ZN(new_n1507_));
  AND3_X1   g1065(.A1(new_n1505_), .A2(new_n1506_), .A3(new_n1507_), .ZN(new_n1508_));
  AOI21_X1  g1066(.A(new_n1506_), .B1(new_n1505_), .B2(new_n1507_), .ZN(new_n1509_));
  OAI21_X1  g1067(.A(new_n1504_), .B1(new_n1508_), .B2(new_n1509_), .ZN(G418));
  NAND2_X1  g1068(.A1(new_n1484_), .A2(new_n811_), .ZN(new_n1511_));
  NAND2_X1  g1069(.A1(new_n1511_), .A2(new_n875_), .ZN(new_n1512_));
  INV_X1    g1070(.A(new_n1512_), .ZN(new_n1513_));
  OAI21_X1  g1071(.A(new_n862_), .B1(new_n1513_), .B2(new_n824_), .ZN(G273));
  OAI21_X1  g1072(.A(new_n857_), .B1(new_n684_), .B2(new_n770_), .ZN(new_n1515_));
  NOR2_X1   g1073(.A1(new_n716_), .A2(new_n702_), .ZN(new_n1516_));
  INV_X1    g1074(.A(new_n827_), .ZN(new_n1517_));
  NAND2_X1  g1075(.A1(new_n1517_), .A2(new_n689_), .ZN(new_n1518_));
  OAI22_X1  g1076(.A1(new_n1516_), .A2(new_n1518_), .B1(new_n688_), .B2(new_n687_), .ZN(new_n1519_));
  NAND2_X1  g1077(.A1(new_n1515_), .A2(new_n1519_), .ZN(new_n1520_));
  OAI21_X1  g1078(.A(new_n1520_), .B1(new_n830_), .B2(new_n1515_), .ZN(new_n1521_));
  INV_X1    g1079(.A(new_n710_), .ZN(new_n1522_));
  XNOR2_X1  g1080(.A(new_n1521_), .B(new_n1522_), .ZN(G298));
  XOR2_X1   g1081(.A(new_n692_), .B(KEYINPUT89), .Z(new_n1524_));
  NOR2_X1   g1082(.A1(new_n1516_), .A2(new_n827_), .ZN(new_n1525_));
  XNOR2_X1  g1083(.A(new_n1524_), .B(new_n1525_), .ZN(new_n1526_));
  NAND2_X1  g1084(.A1(new_n1515_), .A2(new_n1526_), .ZN(new_n1527_));
  NAND2_X1  g1085(.A1(new_n829_), .A2(new_n1517_), .ZN(new_n1528_));
  XOR2_X1   g1086(.A(new_n693_), .B(new_n1528_), .Z(new_n1529_));
  OAI21_X1  g1087(.A(new_n1527_), .B1(new_n1515_), .B2(new_n1529_), .ZN(new_n1530_));
  XOR2_X1   g1088(.A(new_n1530_), .B(KEYINPUT90), .Z(G301));
  INV_X1    g1089(.A(new_n1516_), .ZN(new_n1532_));
  NAND2_X1  g1090(.A1(new_n716_), .A2(new_n702_), .ZN(new_n1533_));
  NAND3_X1  g1091(.A1(new_n1515_), .A2(new_n1532_), .A3(new_n1533_), .ZN(new_n1534_));
  NAND2_X1  g1092(.A1(new_n716_), .A2(new_n698_), .ZN(new_n1535_));
  NAND2_X1  g1093(.A1(new_n1535_), .A2(new_n829_), .ZN(new_n1536_));
  XNOR2_X1  g1094(.A(new_n1536_), .B(KEYINPUT91), .ZN(new_n1537_));
  OAI21_X1  g1095(.A(new_n1534_), .B1(new_n1515_), .B2(new_n1537_), .ZN(G304));
  XNOR2_X1  g1096(.A(new_n1515_), .B(new_n704_), .ZN(G307));
  INV_X1    g1097(.A(new_n680_), .ZN(new_n1540_));
  XNOR2_X1  g1098(.A(new_n678_), .B(new_n1540_), .ZN(G344));
  INV_X1    g1099(.A(G1496), .ZN(new_n1542_));
  MUX2_X1   g1100(.A(new_n1542_), .B(new_n819_), .S(new_n822_), .Z(new_n1543_));
  NAND2_X1  g1101(.A1(new_n1512_), .A2(new_n1543_), .ZN(new_n1544_));
  INV_X1    g1102(.A(new_n816_), .ZN(new_n1545_));
  AOI22_X1  g1103(.A1(new_n1545_), .A2(new_n820_), .B1(new_n861_), .B2(new_n818_), .ZN(new_n1546_));
  XOR2_X1   g1104(.A(new_n1546_), .B(KEYINPUT92), .Z(new_n1547_));
  OAI21_X1  g1105(.A(new_n1544_), .B1(new_n1512_), .B2(new_n1547_), .ZN(G422));
  OAI21_X1  g1106(.A(new_n1544_), .B1(new_n1512_), .B2(new_n1547_), .ZN(G469));
  XNOR2_X1  g1107(.A(new_n1512_), .B(new_n823_), .ZN(G419));
  XNOR2_X1  g1108(.A(new_n1512_), .B(new_n823_), .ZN(G471));
  INV_X1    g1109(.A(new_n579_), .ZN(new_n1552_));
  AOI21_X1  g1110(.A(new_n1552_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n1553_));
  INV_X1    g1111(.A(new_n1553_), .ZN(new_n1554_));
  NOR2_X1   g1112(.A1(new_n1554_), .A2(new_n573_), .ZN(new_n1555_));
  NOR2_X1   g1113(.A1(new_n678_), .A2(new_n1176_), .ZN(new_n1556_));
  INV_X1    g1114(.A(new_n1556_), .ZN(new_n1557_));
  OAI21_X1  g1115(.A(new_n1555_), .B1(new_n1557_), .B2(new_n1183_), .ZN(new_n1558_));
  XNOR2_X1  g1116(.A(new_n1558_), .B(new_n544_), .ZN(G359));
  AOI22_X1  g1117(.A1(new_n1182_), .A2(new_n571_), .B1(new_n548_), .B2(new_n547_), .ZN(new_n1560_));
  INV_X1    g1118(.A(new_n1560_), .ZN(new_n1561_));
  INV_X1    g1119(.A(new_n679_), .ZN(new_n1562_));
  OAI21_X1  g1120(.A(new_n554_), .B1(new_n678_), .B2(new_n1562_), .ZN(new_n1563_));
  NOR2_X1   g1121(.A1(new_n564_), .A2(new_n561_), .ZN(new_n1564_));
  AOI21_X1  g1122(.A(new_n1561_), .B1(new_n1563_), .B2(new_n1564_), .ZN(new_n1565_));
  XNOR2_X1  g1123(.A(new_n1565_), .B(new_n569_), .ZN(G362));
  OR2_X1    g1124(.A1(new_n1556_), .A2(KEYINPUT93), .ZN(new_n1567_));
  NAND2_X1  g1125(.A1(new_n1556_), .A2(KEYINPUT93), .ZN(new_n1568_));
  INV_X1    g1126(.A(new_n571_), .ZN(new_n1569_));
  NAND2_X1  g1127(.A1(new_n562_), .A2(new_n1569_), .ZN(new_n1570_));
  INV_X1    g1128(.A(new_n1570_), .ZN(new_n1571_));
  NAND3_X1  g1129(.A1(new_n1567_), .A2(new_n1568_), .A3(new_n1571_), .ZN(new_n1572_));
  INV_X1    g1130(.A(new_n1182_), .ZN(new_n1573_));
  XNOR2_X1  g1131(.A(new_n1572_), .B(new_n1573_), .ZN(G365));
  XNOR2_X1  g1132(.A(new_n1563_), .B(new_n561_), .ZN(G368));
  NOR2_X1   g1133(.A1(new_n683_), .A2(new_n583_), .ZN(new_n1576_));
  NAND2_X1  g1134(.A1(new_n1576_), .A2(new_n530_), .ZN(new_n1577_));
  NAND2_X1  g1135(.A1(new_n1322_), .A2(new_n585_), .ZN(new_n1578_));
  NAND3_X1  g1136(.A1(new_n520_), .A2(new_n523_), .A3(new_n1578_), .ZN(new_n1579_));
  XNOR2_X1  g1137(.A(new_n1579_), .B(KEYINPUT94), .ZN(new_n1580_));
  AND2_X1   g1138(.A1(new_n1580_), .A2(new_n518_), .ZN(new_n1581_));
  OAI21_X1  g1139(.A(new_n1577_), .B1(new_n1576_), .B2(new_n1581_), .ZN(new_n1582_));
  XNOR2_X1  g1140(.A(new_n1582_), .B(new_n587_), .ZN(G347));
  INV_X1    g1141(.A(new_n529_), .ZN(new_n1584_));
  AOI21_X1  g1142(.A(new_n516_), .B1(new_n523_), .B2(new_n1584_), .ZN(new_n1585_));
  OR2_X1    g1143(.A1(new_n1576_), .A2(new_n586_), .ZN(new_n1586_));
  INV_X1    g1144(.A(new_n589_), .ZN(new_n1587_));
  OAI21_X1  g1145(.A(new_n1585_), .B1(new_n1586_), .B2(new_n1587_), .ZN(new_n1588_));
  XNOR2_X1  g1146(.A(new_n1588_), .B(new_n584_), .ZN(G350));
  NAND2_X1  g1147(.A1(new_n1322_), .A2(G4420), .ZN(new_n1590_));
  INV_X1    g1148(.A(new_n1590_), .ZN(new_n1591_));
  OAI21_X1  g1149(.A(new_n529_), .B1(new_n1576_), .B2(new_n1591_), .ZN(new_n1592_));
  INV_X1    g1150(.A(new_n523_), .ZN(new_n1593_));
  XNOR2_X1  g1151(.A(new_n1592_), .B(new_n1593_), .ZN(G353));
  XOR2_X1   g1152(.A(new_n1576_), .B(new_n586_), .Z(G356));
  INV_X1    g1153(.A(KEYINPUT108), .ZN(new_n1596_));
  NAND2_X1  g1154(.A1(new_n714_), .A2(new_n699_), .ZN(new_n1597_));
  XNOR2_X1  g1155(.A(new_n701_), .B(new_n715_), .ZN(new_n1598_));
  OAI21_X1  g1156(.A(new_n1597_), .B1(new_n1598_), .B2(new_n699_), .ZN(new_n1599_));
  XNOR2_X1  g1157(.A(new_n830_), .B(new_n1599_), .ZN(new_n1600_));
  NAND3_X1  g1158(.A1(new_n1600_), .A2(KEYINPUT104), .A3(new_n716_), .ZN(new_n1601_));
  OR2_X1    g1159(.A1(new_n830_), .A2(new_n1599_), .ZN(new_n1602_));
  INV_X1    g1160(.A(new_n716_), .ZN(new_n1603_));
  NAND2_X1  g1161(.A1(new_n830_), .A2(new_n1599_), .ZN(new_n1604_));
  NAND3_X1  g1162(.A1(new_n1602_), .A2(new_n1603_), .A3(new_n1604_), .ZN(new_n1605_));
  NAND3_X1  g1163(.A1(new_n1601_), .A2(new_n1522_), .A3(new_n1605_), .ZN(new_n1606_));
  AOI21_X1  g1164(.A(KEYINPUT104), .B1(new_n1600_), .B2(new_n716_), .ZN(new_n1607_));
  OAI21_X1  g1165(.A(KEYINPUT105), .B1(new_n1606_), .B2(new_n1607_), .ZN(new_n1608_));
  INV_X1    g1166(.A(new_n1607_), .ZN(new_n1609_));
  AND2_X1   g1167(.A1(new_n1605_), .A2(new_n1522_), .ZN(new_n1610_));
  INV_X1    g1168(.A(KEYINPUT105), .ZN(new_n1611_));
  NAND4_X1  g1169(.A1(new_n1609_), .A2(new_n1610_), .A3(new_n1611_), .A4(new_n1601_), .ZN(new_n1612_));
  NAND2_X1  g1170(.A1(new_n1600_), .A2(new_n716_), .ZN(new_n1613_));
  AOI21_X1  g1171(.A(new_n1522_), .B1(new_n1613_), .B2(new_n1605_), .ZN(new_n1614_));
  INV_X1    g1172(.A(new_n1614_), .ZN(new_n1615_));
  NAND3_X1  g1173(.A1(new_n1608_), .A2(new_n1612_), .A3(new_n1615_), .ZN(new_n1616_));
  INV_X1    g1174(.A(new_n692_), .ZN(new_n1617_));
  INV_X1    g1175(.A(KEYINPUT106), .ZN(new_n1618_));
  NAND2_X1  g1176(.A1(new_n1617_), .A2(new_n1618_), .ZN(new_n1619_));
  NAND2_X1  g1177(.A1(new_n692_), .A2(KEYINPUT106), .ZN(new_n1620_));
  NAND3_X1  g1178(.A1(new_n1616_), .A2(new_n1619_), .A3(new_n1620_), .ZN(new_n1621_));
  NAND3_X1  g1179(.A1(new_n1609_), .A2(new_n1610_), .A3(new_n1601_), .ZN(new_n1622_));
  AOI21_X1  g1180(.A(new_n1614_), .B1(new_n1622_), .B2(KEYINPUT105), .ZN(new_n1623_));
  NAND4_X1  g1181(.A1(new_n1623_), .A2(new_n1618_), .A3(new_n1617_), .A4(new_n1612_), .ZN(new_n1624_));
  NOR2_X1   g1182(.A1(new_n856_), .A2(new_n769_), .ZN(new_n1625_));
  NAND3_X1  g1183(.A1(new_n1621_), .A2(new_n1624_), .A3(new_n1625_), .ZN(new_n1626_));
  NAND2_X1  g1184(.A1(new_n1617_), .A2(KEYINPUT102), .ZN(new_n1627_));
  XNOR2_X1  g1185(.A(new_n1519_), .B(new_n1522_), .ZN(new_n1628_));
  AOI21_X1  g1186(.A(new_n702_), .B1(new_n713_), .B2(G2247), .ZN(new_n1629_));
  AND2_X1   g1187(.A1(new_n702_), .A2(new_n715_), .ZN(new_n1630_));
  OAI21_X1  g1188(.A(new_n716_), .B1(new_n1629_), .B2(new_n1630_), .ZN(new_n1631_));
  XNOR2_X1  g1189(.A(new_n1631_), .B(new_n703_), .ZN(new_n1632_));
  NOR2_X1   g1190(.A1(new_n1628_), .A2(new_n1632_), .ZN(new_n1633_));
  OR2_X1    g1191(.A1(new_n1519_), .A2(new_n710_), .ZN(new_n1634_));
  NAND2_X1  g1192(.A1(new_n1519_), .A2(new_n710_), .ZN(new_n1635_));
  AND3_X1   g1193(.A1(new_n1634_), .A2(new_n1632_), .A3(new_n1635_), .ZN(new_n1636_));
  OAI21_X1  g1194(.A(new_n1627_), .B1(new_n1633_), .B2(new_n1636_), .ZN(new_n1637_));
  NAND2_X1  g1195(.A1(new_n1634_), .A2(new_n1635_), .ZN(new_n1638_));
  INV_X1    g1196(.A(new_n1632_), .ZN(new_n1639_));
  NAND2_X1  g1197(.A1(new_n1638_), .A2(new_n1639_), .ZN(new_n1640_));
  NAND2_X1  g1198(.A1(new_n1628_), .A2(new_n1632_), .ZN(new_n1641_));
  XOR2_X1   g1199(.A(new_n692_), .B(KEYINPUT102), .Z(new_n1642_));
  NAND3_X1  g1200(.A1(new_n1640_), .A2(new_n1641_), .A3(new_n1642_), .ZN(new_n1643_));
  NAND2_X1  g1201(.A1(new_n1637_), .A2(new_n1643_), .ZN(new_n1644_));
  OAI21_X1  g1202(.A(new_n1644_), .B1(new_n769_), .B2(new_n856_), .ZN(new_n1645_));
  NAND2_X1  g1203(.A1(new_n1626_), .A2(new_n1645_), .ZN(new_n1646_));
  NAND2_X1  g1204(.A1(new_n1198_), .A2(new_n1194_), .ZN(new_n1647_));
  INV_X1    g1205(.A(new_n1193_), .ZN(new_n1648_));
  NAND2_X1  g1206(.A1(new_n1647_), .A2(new_n1648_), .ZN(new_n1649_));
  NAND2_X1  g1207(.A1(new_n1646_), .A2(new_n1649_), .ZN(new_n1650_));
  AND2_X1   g1208(.A1(new_n1621_), .A2(new_n1624_), .ZN(new_n1651_));
  NOR2_X1   g1209(.A1(new_n1649_), .A2(new_n856_), .ZN(new_n1652_));
  AOI21_X1  g1210(.A(new_n857_), .B1(new_n1637_), .B2(new_n1643_), .ZN(new_n1653_));
  NAND3_X1  g1211(.A1(new_n1647_), .A2(new_n1653_), .A3(new_n1648_), .ZN(new_n1654_));
  NAND2_X1  g1212(.A1(new_n1654_), .A2(KEYINPUT103), .ZN(new_n1655_));
  INV_X1    g1213(.A(KEYINPUT103), .ZN(new_n1656_));
  NAND3_X1  g1214(.A1(new_n1199_), .A2(new_n1656_), .A3(new_n1653_), .ZN(new_n1657_));
  AOI22_X1  g1215(.A1(new_n1651_), .A2(new_n1652_), .B1(new_n1655_), .B2(new_n1657_), .ZN(new_n1658_));
  INV_X1    g1216(.A(KEYINPUT107), .ZN(new_n1659_));
  NAND3_X1  g1217(.A1(new_n1650_), .A2(new_n1658_), .A3(new_n1659_), .ZN(new_n1660_));
  NAND2_X1  g1218(.A1(new_n1655_), .A2(new_n1657_), .ZN(new_n1661_));
  NAND4_X1  g1219(.A1(new_n1621_), .A2(new_n1624_), .A3(new_n1199_), .A4(new_n857_), .ZN(new_n1662_));
  NAND2_X1  g1220(.A1(new_n1661_), .A2(new_n1662_), .ZN(new_n1663_));
  AOI21_X1  g1221(.A(new_n1199_), .B1(new_n1626_), .B2(new_n1645_), .ZN(new_n1664_));
  OAI21_X1  g1222(.A(KEYINPUT107), .B1(new_n1663_), .B2(new_n1664_), .ZN(new_n1665_));
  AND2_X1   g1223(.A1(new_n1660_), .A2(new_n1665_), .ZN(new_n1666_));
  OAI21_X1  g1224(.A(new_n841_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n1667_));
  NAND3_X1  g1225(.A1(new_n749_), .A2(G2211), .A3(new_n742_), .ZN(new_n1668_));
  NAND3_X1  g1226(.A1(new_n1478_), .A2(new_n839_), .A3(new_n1668_), .ZN(new_n1669_));
  OAI22_X1  g1227(.A1(new_n1667_), .A2(new_n1669_), .B1(new_n848_), .B2(new_n842_), .ZN(new_n1670_));
  OAI211_X1 g1228(.A(new_n835_), .B(new_n841_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n1671_));
  INV_X1    g1229(.A(new_n854_), .ZN(new_n1672_));
  NAND2_X1  g1230(.A1(new_n1671_), .A2(new_n1672_), .ZN(new_n1673_));
  NOR2_X1   g1231(.A1(new_n1670_), .A2(new_n1673_), .ZN(new_n1674_));
  AOI21_X1  g1232(.A(new_n1458_), .B1(new_n1674_), .B2(KEYINPUT95), .ZN(new_n1675_));
  INV_X1    g1233(.A(KEYINPUT95), .ZN(new_n1676_));
  OAI21_X1  g1234(.A(new_n1676_), .B1(new_n1670_), .B2(new_n1673_), .ZN(new_n1677_));
  OAI21_X1  g1235(.A(new_n1668_), .B1(new_n725_), .B2(new_n758_), .ZN(new_n1678_));
  NAND2_X1  g1236(.A1(new_n836_), .A2(new_n1678_), .ZN(new_n1679_));
  NOR3_X1   g1237(.A1(new_n832_), .A2(new_n834_), .A3(new_n840_), .ZN(new_n1680_));
  OAI21_X1  g1238(.A(new_n1668_), .B1(new_n1680_), .B2(new_n721_), .ZN(new_n1681_));
  NAND2_X1  g1239(.A1(new_n1679_), .A2(new_n1681_), .ZN(new_n1682_));
  NOR2_X1   g1240(.A1(new_n1479_), .A2(new_n759_), .ZN(new_n1683_));
  NAND2_X1  g1241(.A1(new_n1682_), .A2(new_n1683_), .ZN(new_n1684_));
  OAI211_X1 g1242(.A(new_n1679_), .B(new_n1681_), .C1(new_n759_), .C2(new_n1479_), .ZN(new_n1685_));
  AOI22_X1  g1243(.A1(new_n1675_), .A2(new_n1677_), .B1(new_n1684_), .B2(new_n1685_), .ZN(new_n1686_));
  NAND4_X1  g1244(.A1(new_n1460_), .A2(KEYINPUT95), .A3(new_n760_), .A4(new_n1462_), .ZN(new_n1687_));
  NAND3_X1  g1245(.A1(new_n1677_), .A2(new_n1687_), .A3(new_n1459_), .ZN(new_n1688_));
  NAND2_X1  g1246(.A1(new_n1684_), .A2(new_n1685_), .ZN(new_n1689_));
  NOR2_X1   g1247(.A1(new_n1688_), .A2(new_n1689_), .ZN(new_n1690_));
  OAI21_X1  g1248(.A(new_n1446_), .B1(new_n1686_), .B2(new_n1690_), .ZN(new_n1691_));
  NAND4_X1  g1249(.A1(new_n1675_), .A2(new_n1677_), .A3(new_n1684_), .A4(new_n1685_), .ZN(new_n1692_));
  NAND2_X1  g1250(.A1(new_n1688_), .A2(new_n1689_), .ZN(new_n1693_));
  NAND3_X1  g1251(.A1(new_n1692_), .A2(new_n1465_), .A3(new_n1693_), .ZN(new_n1694_));
  NAND3_X1  g1252(.A1(new_n1691_), .A2(KEYINPUT96), .A3(new_n1694_), .ZN(new_n1695_));
  INV_X1    g1253(.A(KEYINPUT96), .ZN(new_n1696_));
  NAND4_X1  g1254(.A1(new_n1692_), .A2(new_n1696_), .A3(new_n1693_), .A4(new_n1465_), .ZN(new_n1697_));
  NAND3_X1  g1255(.A1(new_n1695_), .A2(new_n839_), .A3(new_n1697_), .ZN(new_n1698_));
  AND2_X1   g1256(.A1(new_n1698_), .A2(new_n768_), .ZN(new_n1699_));
  INV_X1    g1257(.A(KEYINPUT97), .ZN(new_n1700_));
  NAND3_X1  g1258(.A1(new_n1691_), .A2(new_n1700_), .A3(new_n1694_), .ZN(new_n1701_));
  OAI211_X1 g1259(.A(KEYINPUT97), .B(new_n1446_), .C1(new_n1686_), .C2(new_n1690_), .ZN(new_n1702_));
  NAND2_X1  g1260(.A1(new_n1701_), .A2(new_n1702_), .ZN(new_n1703_));
  NAND2_X1  g1261(.A1(new_n1703_), .A2(new_n758_), .ZN(new_n1704_));
  AOI21_X1  g1262(.A(new_n725_), .B1(new_n1699_), .B2(new_n1704_), .ZN(new_n1705_));
  AND3_X1   g1263(.A1(new_n1701_), .A2(new_n839_), .A3(new_n1702_), .ZN(new_n1706_));
  AOI21_X1  g1264(.A(new_n839_), .B1(new_n1695_), .B2(new_n1697_), .ZN(new_n1707_));
  OAI21_X1  g1265(.A(new_n767_), .B1(new_n1706_), .B2(new_n1707_), .ZN(new_n1708_));
  INV_X1    g1266(.A(KEYINPUT98), .ZN(new_n1709_));
  NAND2_X1  g1267(.A1(new_n1708_), .A2(new_n1709_), .ZN(new_n1710_));
  OAI211_X1 g1268(.A(KEYINPUT98), .B(new_n767_), .C1(new_n1706_), .C2(new_n1707_), .ZN(new_n1711_));
  NAND3_X1  g1269(.A1(new_n1705_), .A2(new_n1710_), .A3(new_n1711_), .ZN(new_n1712_));
  NAND2_X1  g1270(.A1(new_n1695_), .A2(new_n1697_), .ZN(new_n1713_));
  NAND2_X1  g1271(.A1(new_n1713_), .A2(new_n758_), .ZN(new_n1714_));
  NAND3_X1  g1272(.A1(new_n1701_), .A2(new_n839_), .A3(new_n1702_), .ZN(new_n1715_));
  NAND3_X1  g1273(.A1(new_n1714_), .A2(new_n768_), .A3(new_n1715_), .ZN(new_n1716_));
  NAND2_X1  g1274(.A1(new_n1708_), .A2(new_n1716_), .ZN(new_n1717_));
  NAND2_X1  g1275(.A1(new_n1717_), .A2(new_n725_), .ZN(new_n1718_));
  AND3_X1   g1276(.A1(new_n1712_), .A2(new_n1461_), .A3(new_n1718_), .ZN(new_n1719_));
  AOI21_X1  g1277(.A(new_n1461_), .B1(new_n1712_), .B2(new_n1718_), .ZN(new_n1720_));
  OAI21_X1  g1278(.A(new_n1649_), .B1(new_n1719_), .B2(new_n1720_), .ZN(new_n1721_));
  XNOR2_X1  g1279(.A(new_n1479_), .B(new_n758_), .ZN(new_n1722_));
  NAND2_X1  g1280(.A1(new_n843_), .A2(new_n750_), .ZN(new_n1723_));
  INV_X1    g1281(.A(KEYINPUT99), .ZN(new_n1724_));
  AOI21_X1  g1282(.A(new_n1724_), .B1(new_n836_), .B2(new_n1478_), .ZN(new_n1725_));
  NAND2_X1  g1283(.A1(new_n1723_), .A2(new_n1725_), .ZN(new_n1726_));
  NAND3_X1  g1284(.A1(new_n843_), .A2(new_n1724_), .A3(new_n750_), .ZN(new_n1727_));
  NAND3_X1  g1285(.A1(new_n1722_), .A2(new_n1726_), .A3(new_n1727_), .ZN(new_n1728_));
  INV_X1    g1286(.A(new_n1728_), .ZN(new_n1729_));
  AOI21_X1  g1287(.A(new_n1722_), .B1(new_n1726_), .B2(new_n1727_), .ZN(new_n1730_));
  OAI21_X1  g1288(.A(new_n1446_), .B1(new_n1729_), .B2(new_n1730_), .ZN(new_n1731_));
  NAND2_X1  g1289(.A1(new_n1726_), .A2(new_n1727_), .ZN(new_n1732_));
  INV_X1    g1290(.A(new_n1722_), .ZN(new_n1733_));
  NAND2_X1  g1291(.A1(new_n1732_), .A2(new_n1733_), .ZN(new_n1734_));
  NAND3_X1  g1292(.A1(new_n1734_), .A2(new_n1465_), .A3(new_n1728_), .ZN(new_n1735_));
  NAND3_X1  g1293(.A1(new_n1731_), .A2(new_n1464_), .A3(new_n1735_), .ZN(new_n1736_));
  INV_X1    g1294(.A(new_n1736_), .ZN(new_n1737_));
  AOI21_X1  g1295(.A(new_n1464_), .B1(new_n1731_), .B2(new_n1735_), .ZN(new_n1738_));
  OAI21_X1  g1296(.A(new_n767_), .B1(new_n1737_), .B2(new_n1738_), .ZN(new_n1739_));
  INV_X1    g1297(.A(KEYINPUT100), .ZN(new_n1740_));
  NAND2_X1  g1298(.A1(new_n1731_), .A2(new_n1735_), .ZN(new_n1741_));
  NAND2_X1  g1299(.A1(new_n1741_), .A2(new_n1463_), .ZN(new_n1742_));
  NAND3_X1  g1300(.A1(new_n1742_), .A2(new_n768_), .A3(new_n1736_), .ZN(new_n1743_));
  NAND3_X1  g1301(.A1(new_n1739_), .A2(new_n1740_), .A3(new_n1743_), .ZN(new_n1744_));
  NAND4_X1  g1302(.A1(new_n1742_), .A2(KEYINPUT100), .A3(new_n1736_), .A4(new_n768_), .ZN(new_n1745_));
  NAND3_X1  g1303(.A1(new_n1744_), .A2(new_n725_), .A3(new_n1745_), .ZN(new_n1746_));
  NAND4_X1  g1304(.A1(new_n1739_), .A2(new_n1743_), .A3(KEYINPUT101), .A4(new_n841_), .ZN(new_n1747_));
  NAND3_X1  g1305(.A1(new_n1739_), .A2(new_n841_), .A3(new_n1743_), .ZN(new_n1748_));
  INV_X1    g1306(.A(KEYINPUT101), .ZN(new_n1749_));
  NAND2_X1  g1307(.A1(new_n1748_), .A2(new_n1749_), .ZN(new_n1750_));
  NAND3_X1  g1308(.A1(new_n1746_), .A2(new_n1747_), .A3(new_n1750_), .ZN(new_n1751_));
  NAND2_X1  g1309(.A1(new_n1751_), .A2(new_n848_), .ZN(new_n1752_));
  NAND4_X1  g1310(.A1(new_n1746_), .A2(new_n1750_), .A3(new_n1461_), .A4(new_n1747_), .ZN(new_n1753_));
  NAND3_X1  g1311(.A1(new_n1752_), .A2(new_n1199_), .A3(new_n1753_), .ZN(new_n1754_));
  AOI21_X1  g1312(.A(new_n1666_), .B1(new_n1721_), .B2(new_n1754_), .ZN(new_n1755_));
  NAND2_X1  g1313(.A1(new_n1650_), .A2(new_n1658_), .ZN(new_n1756_));
  NAND2_X1  g1314(.A1(new_n1754_), .A2(new_n1756_), .ZN(new_n1757_));
  NAND3_X1  g1315(.A1(new_n1712_), .A2(new_n1461_), .A3(new_n1718_), .ZN(new_n1758_));
  AOI21_X1  g1316(.A(new_n1461_), .B1(new_n1717_), .B2(new_n841_), .ZN(new_n1759_));
  AOI21_X1  g1317(.A(new_n841_), .B1(new_n1699_), .B2(new_n1704_), .ZN(new_n1760_));
  NAND3_X1  g1318(.A1(new_n1760_), .A2(new_n1710_), .A3(new_n1711_), .ZN(new_n1761_));
  NAND2_X1  g1319(.A1(new_n1759_), .A2(new_n1761_), .ZN(new_n1762_));
  NAND2_X1  g1320(.A1(new_n1758_), .A2(new_n1762_), .ZN(new_n1763_));
  AOI21_X1  g1321(.A(new_n1757_), .B1(new_n1649_), .B2(new_n1763_), .ZN(new_n1764_));
  OAI21_X1  g1322(.A(new_n1596_), .B1(new_n1755_), .B2(new_n1764_), .ZN(new_n1765_));
  NAND2_X1  g1323(.A1(new_n1763_), .A2(new_n1649_), .ZN(new_n1766_));
  NAND3_X1  g1324(.A1(new_n1766_), .A2(new_n1754_), .A3(new_n1756_), .ZN(new_n1767_));
  INV_X1    g1325(.A(new_n1754_), .ZN(new_n1768_));
  NAND2_X1  g1326(.A1(new_n1712_), .A2(new_n1718_), .ZN(new_n1769_));
  NAND2_X1  g1327(.A1(new_n1769_), .A2(new_n848_), .ZN(new_n1770_));
  NAND2_X1  g1328(.A1(new_n1770_), .A2(new_n1758_), .ZN(new_n1771_));
  AOI21_X1  g1329(.A(new_n1768_), .B1(new_n1771_), .B2(new_n1649_), .ZN(new_n1772_));
  OAI211_X1 g1330(.A(KEYINPUT108), .B(new_n1767_), .C1(new_n1772_), .C2(new_n1666_), .ZN(new_n1773_));
  NAND2_X1  g1331(.A1(new_n1765_), .A2(new_n1773_), .ZN(G321));
  INV_X1    g1332(.A(new_n1455_), .ZN(new_n1775_));
  INV_X1    g1333(.A(KEYINPUT109), .ZN(new_n1776_));
  NAND2_X1  g1334(.A1(new_n868_), .A2(new_n1776_), .ZN(new_n1777_));
  NAND2_X1  g1335(.A1(new_n803_), .A2(new_n796_), .ZN(new_n1778_));
  NAND3_X1  g1336(.A1(new_n863_), .A2(KEYINPUT109), .A3(new_n867_), .ZN(new_n1779_));
  AND3_X1   g1337(.A1(new_n1777_), .A2(new_n1778_), .A3(new_n1779_), .ZN(new_n1780_));
  NAND3_X1  g1338(.A1(new_n787_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n1781_));
  NAND2_X1  g1339(.A1(new_n1781_), .A2(new_n871_), .ZN(new_n1782_));
  NAND2_X1  g1340(.A1(new_n1782_), .A2(new_n802_), .ZN(new_n1783_));
  INV_X1    g1341(.A(new_n802_), .ZN(new_n1784_));
  NAND4_X1  g1342(.A1(new_n1494_), .A2(new_n1781_), .A3(new_n1784_), .A4(new_n871_), .ZN(new_n1785_));
  NAND2_X1  g1343(.A1(new_n1783_), .A2(new_n1785_), .ZN(new_n1786_));
  NAND3_X1  g1344(.A1(new_n1780_), .A2(KEYINPUT110), .A3(new_n1786_), .ZN(new_n1787_));
  INV_X1    g1345(.A(new_n1786_), .ZN(new_n1788_));
  NAND4_X1  g1346(.A1(new_n1777_), .A2(KEYINPUT110), .A3(new_n1778_), .A4(new_n1779_), .ZN(new_n1789_));
  NAND2_X1  g1347(.A1(new_n1788_), .A2(new_n1789_), .ZN(new_n1790_));
  NAND2_X1  g1348(.A1(new_n1787_), .A2(new_n1790_), .ZN(new_n1791_));
  NAND2_X1  g1349(.A1(new_n1488_), .A2(new_n804_), .ZN(new_n1792_));
  NAND2_X1  g1350(.A1(new_n1791_), .A2(new_n1792_), .ZN(new_n1793_));
  INV_X1    g1351(.A(new_n1792_), .ZN(new_n1794_));
  INV_X1    g1352(.A(new_n1779_), .ZN(new_n1795_));
  AOI21_X1  g1353(.A(KEYINPUT109), .B1(new_n863_), .B2(new_n867_), .ZN(new_n1796_));
  NOR2_X1   g1354(.A1(new_n1795_), .A2(new_n1796_), .ZN(new_n1797_));
  NAND2_X1  g1355(.A1(new_n1797_), .A2(new_n1778_), .ZN(new_n1798_));
  NAND2_X1  g1356(.A1(new_n1798_), .A2(new_n1788_), .ZN(new_n1799_));
  NAND2_X1  g1357(.A1(new_n1780_), .A2(new_n1786_), .ZN(new_n1800_));
  NAND3_X1  g1358(.A1(new_n1794_), .A2(new_n1799_), .A3(new_n1800_), .ZN(new_n1801_));
  NAND3_X1  g1359(.A1(new_n1793_), .A2(new_n803_), .A3(new_n1801_), .ZN(new_n1802_));
  NAND3_X1  g1360(.A1(new_n1799_), .A2(new_n1800_), .A3(new_n1792_), .ZN(new_n1803_));
  INV_X1    g1361(.A(new_n803_), .ZN(new_n1804_));
  XNOR2_X1  g1362(.A(new_n1789_), .B(new_n1786_), .ZN(new_n1805_));
  OAI211_X1 g1363(.A(new_n1803_), .B(new_n1804_), .C1(new_n1805_), .C2(new_n1792_), .ZN(new_n1806_));
  NAND3_X1  g1364(.A1(new_n1802_), .A2(new_n1806_), .A3(new_n796_), .ZN(new_n1807_));
  INV_X1    g1365(.A(new_n1807_), .ZN(new_n1808_));
  AND3_X1   g1366(.A1(new_n1794_), .A2(new_n1799_), .A3(new_n1800_), .ZN(new_n1809_));
  AOI21_X1  g1367(.A(new_n1794_), .B1(new_n1787_), .B2(new_n1790_), .ZN(new_n1810_));
  OAI21_X1  g1368(.A(new_n1804_), .B1(new_n1809_), .B2(new_n1810_), .ZN(new_n1811_));
  AOI21_X1  g1369(.A(new_n796_), .B1(new_n1811_), .B2(new_n1802_), .ZN(new_n1812_));
  NOR3_X1   g1370(.A1(new_n1808_), .A2(new_n1812_), .A3(new_n812_), .ZN(new_n1813_));
  INV_X1    g1371(.A(new_n1802_), .ZN(new_n1814_));
  AOI21_X1  g1372(.A(new_n803_), .B1(new_n1793_), .B2(new_n1801_), .ZN(new_n1815_));
  OAI21_X1  g1373(.A(new_n795_), .B1(new_n1814_), .B2(new_n1815_), .ZN(new_n1816_));
  AOI21_X1  g1374(.A(new_n811_), .B1(new_n1816_), .B2(new_n1807_), .ZN(new_n1817_));
  OAI21_X1  g1375(.A(new_n788_), .B1(new_n1813_), .B2(new_n1817_), .ZN(new_n1818_));
  NAND2_X1  g1376(.A1(new_n1818_), .A2(KEYINPUT111), .ZN(new_n1819_));
  OAI21_X1  g1377(.A(new_n812_), .B1(new_n1808_), .B2(new_n1812_), .ZN(new_n1820_));
  NAND3_X1  g1378(.A1(new_n1816_), .A2(new_n811_), .A3(new_n1807_), .ZN(new_n1821_));
  NAND2_X1  g1379(.A1(new_n1820_), .A2(new_n1821_), .ZN(new_n1822_));
  INV_X1    g1380(.A(KEYINPUT111), .ZN(new_n1823_));
  NAND3_X1  g1381(.A1(new_n1822_), .A2(new_n1823_), .A3(new_n788_), .ZN(new_n1824_));
  NAND2_X1  g1382(.A1(new_n1819_), .A2(new_n1824_), .ZN(new_n1825_));
  OAI21_X1  g1383(.A(new_n796_), .B1(new_n1814_), .B2(new_n1815_), .ZN(new_n1826_));
  NAND3_X1  g1384(.A1(new_n1802_), .A2(new_n1806_), .A3(new_n795_), .ZN(new_n1827_));
  NAND3_X1  g1385(.A1(new_n1826_), .A2(new_n812_), .A3(new_n1827_), .ZN(new_n1828_));
  NAND3_X1  g1386(.A1(new_n1821_), .A2(new_n1828_), .A3(new_n787_), .ZN(new_n1829_));
  NAND2_X1  g1387(.A1(new_n1829_), .A2(KEYINPUT112), .ZN(new_n1830_));
  INV_X1    g1388(.A(KEYINPUT112), .ZN(new_n1831_));
  NAND4_X1  g1389(.A1(new_n1821_), .A2(new_n1828_), .A3(new_n1831_), .A4(new_n787_), .ZN(new_n1832_));
  NAND2_X1  g1390(.A1(new_n1830_), .A2(new_n1832_), .ZN(new_n1833_));
  NAND3_X1  g1391(.A1(new_n1825_), .A2(new_n778_), .A3(new_n1833_), .ZN(new_n1834_));
  NAND2_X1  g1392(.A1(new_n1822_), .A2(new_n787_), .ZN(new_n1835_));
  NAND3_X1  g1393(.A1(new_n1821_), .A2(new_n1828_), .A3(new_n788_), .ZN(new_n1836_));
  NAND3_X1  g1394(.A1(new_n1835_), .A2(new_n779_), .A3(new_n1836_), .ZN(new_n1837_));
  AOI21_X1  g1395(.A(new_n1775_), .B1(new_n1834_), .B2(new_n1837_), .ZN(new_n1838_));
  INV_X1    g1396(.A(new_n1494_), .ZN(new_n1839_));
  OAI21_X1  g1397(.A(new_n1485_), .B1(new_n1782_), .B2(new_n1839_), .ZN(new_n1840_));
  NAND3_X1  g1398(.A1(new_n1781_), .A2(new_n800_), .A3(new_n871_), .ZN(new_n1841_));
  NAND3_X1  g1399(.A1(new_n1797_), .A2(new_n1840_), .A3(new_n1841_), .ZN(new_n1842_));
  INV_X1    g1400(.A(new_n1842_), .ZN(new_n1843_));
  AOI21_X1  g1401(.A(new_n1797_), .B1(new_n1840_), .B2(new_n1841_), .ZN(new_n1844_));
  OAI21_X1  g1402(.A(new_n1489_), .B1(new_n1843_), .B2(new_n1844_), .ZN(new_n1845_));
  NAND2_X1  g1403(.A1(new_n1840_), .A2(new_n1841_), .ZN(new_n1846_));
  NAND2_X1  g1404(.A1(new_n1486_), .A2(new_n793_), .ZN(new_n1847_));
  NAND2_X1  g1405(.A1(new_n1846_), .A2(new_n1847_), .ZN(new_n1848_));
  NAND3_X1  g1406(.A1(new_n1842_), .A2(new_n1848_), .A3(new_n1488_), .ZN(new_n1849_));
  AND3_X1   g1407(.A1(new_n1845_), .A2(new_n803_), .A3(new_n1849_), .ZN(new_n1850_));
  AOI21_X1  g1408(.A(new_n803_), .B1(new_n1845_), .B2(new_n1849_), .ZN(new_n1851_));
  OAI21_X1  g1409(.A(new_n796_), .B1(new_n1850_), .B2(new_n1851_), .ZN(new_n1852_));
  NAND3_X1  g1410(.A1(new_n1845_), .A2(new_n803_), .A3(new_n1849_), .ZN(new_n1853_));
  OAI21_X1  g1411(.A(new_n1488_), .B1(new_n1843_), .B2(new_n1844_), .ZN(new_n1854_));
  NAND3_X1  g1412(.A1(new_n1842_), .A2(new_n1848_), .A3(new_n1489_), .ZN(new_n1855_));
  NAND3_X1  g1413(.A1(new_n1854_), .A2(new_n1804_), .A3(new_n1855_), .ZN(new_n1856_));
  NAND3_X1  g1414(.A1(new_n1853_), .A2(new_n1856_), .A3(new_n795_), .ZN(new_n1857_));
  AND4_X1   g1415(.A1(new_n812_), .A2(new_n1852_), .A3(new_n787_), .A4(new_n1857_), .ZN(new_n1858_));
  OAI21_X1  g1416(.A(new_n795_), .B1(new_n1850_), .B2(new_n1851_), .ZN(new_n1859_));
  NAND3_X1  g1417(.A1(new_n1853_), .A2(new_n1856_), .A3(new_n796_), .ZN(new_n1860_));
  NAND3_X1  g1418(.A1(new_n1859_), .A2(new_n811_), .A3(new_n1860_), .ZN(new_n1861_));
  AOI21_X1  g1419(.A(new_n811_), .B1(new_n1859_), .B2(new_n1860_), .ZN(new_n1862_));
  NAND2_X1  g1420(.A1(new_n788_), .A2(KEYINPUT113), .ZN(new_n1863_));
  OAI21_X1  g1421(.A(new_n1861_), .B1(new_n1862_), .B2(new_n1863_), .ZN(new_n1864_));
  INV_X1    g1422(.A(new_n1863_), .ZN(new_n1865_));
  NAND4_X1  g1423(.A1(new_n1859_), .A2(new_n811_), .A3(new_n1860_), .A4(new_n1865_), .ZN(new_n1866_));
  AOI21_X1  g1424(.A(new_n1858_), .B1(new_n1864_), .B2(new_n1866_), .ZN(new_n1867_));
  NOR2_X1   g1425(.A1(new_n1867_), .A2(new_n778_), .ZN(new_n1868_));
  AOI211_X1 g1426(.A(new_n779_), .B(new_n1858_), .C1(new_n1864_), .C2(new_n1866_), .ZN(new_n1869_));
  OAI21_X1  g1427(.A(new_n1775_), .B1(new_n1868_), .B2(new_n1869_), .ZN(new_n1870_));
  AND2_X1   g1428(.A1(new_n875_), .A2(new_n1543_), .ZN(new_n1871_));
  NAND2_X1  g1429(.A1(new_n1775_), .A2(new_n1871_), .ZN(new_n1872_));
  XNOR2_X1  g1430(.A(new_n1872_), .B(KEYINPUT114), .ZN(new_n1873_));
  NAND2_X1  g1431(.A1(new_n874_), .A2(new_n1546_), .ZN(new_n1874_));
  NAND2_X1  g1432(.A1(new_n814_), .A2(new_n875_), .ZN(new_n1875_));
  AOI22_X1  g1433(.A1(new_n1871_), .A2(new_n814_), .B1(new_n1875_), .B2(new_n1546_), .ZN(new_n1876_));
  MUX2_X1   g1434(.A(new_n1874_), .B(new_n1876_), .S(new_n1455_), .Z(new_n1877_));
  NAND2_X1  g1435(.A1(new_n1873_), .A2(new_n1877_), .ZN(new_n1878_));
  NAND2_X1  g1436(.A1(new_n1870_), .A2(new_n1878_), .ZN(new_n1879_));
  NOR2_X1   g1437(.A1(new_n1838_), .A2(new_n1879_), .ZN(new_n1880_));
  AND3_X1   g1438(.A1(new_n1825_), .A2(new_n778_), .A3(new_n1833_), .ZN(new_n1881_));
  AOI21_X1  g1439(.A(new_n778_), .B1(new_n1825_), .B2(new_n1833_), .ZN(new_n1882_));
  OAI21_X1  g1440(.A(new_n1455_), .B1(new_n1881_), .B2(new_n1882_), .ZN(new_n1883_));
  NAND2_X1  g1441(.A1(new_n1883_), .A2(new_n1870_), .ZN(new_n1884_));
  INV_X1    g1442(.A(new_n1878_), .ZN(new_n1885_));
  AOI21_X1  g1443(.A(new_n1880_), .B1(new_n1884_), .B2(new_n1885_), .ZN(G338));
  INV_X1    g1444(.A(new_n1174_), .ZN(new_n1887_));
  OAI21_X1  g1445(.A(new_n665_), .B1(new_n505_), .B2(new_n1887_), .ZN(new_n1888_));
  AOI21_X1  g1446(.A(new_n622_), .B1(new_n1186_), .B2(new_n1888_), .ZN(new_n1889_));
  INV_X1    g1447(.A(new_n1889_), .ZN(new_n1890_));
  NAND3_X1  g1448(.A1(new_n1553_), .A2(new_n682_), .A3(new_n572_), .ZN(new_n1891_));
  NAND2_X1  g1449(.A1(new_n1891_), .A2(KEYINPUT115), .ZN(new_n1892_));
  INV_X1    g1450(.A(KEYINPUT115), .ZN(new_n1893_));
  NAND4_X1  g1451(.A1(new_n1553_), .A2(new_n1893_), .A3(new_n682_), .A4(new_n572_), .ZN(new_n1894_));
  NOR2_X1   g1452(.A1(new_n1560_), .A2(new_n1562_), .ZN(new_n1895_));
  INV_X1    g1453(.A(new_n1895_), .ZN(new_n1896_));
  OAI21_X1  g1454(.A(new_n679_), .B1(new_n564_), .B2(new_n561_), .ZN(new_n1897_));
  NAND2_X1  g1455(.A1(new_n1560_), .A2(new_n1897_), .ZN(new_n1898_));
  NAND2_X1  g1456(.A1(new_n1571_), .A2(new_n1176_), .ZN(new_n1899_));
  NAND3_X1  g1457(.A1(new_n1896_), .A2(new_n1898_), .A3(new_n1899_), .ZN(new_n1900_));
  INV_X1    g1458(.A(new_n1900_), .ZN(new_n1901_));
  AOI21_X1  g1459(.A(new_n1899_), .B1(new_n1896_), .B2(new_n1898_), .ZN(new_n1902_));
  OAI211_X1 g1460(.A(new_n1892_), .B(new_n1894_), .C1(new_n1901_), .C2(new_n1902_), .ZN(new_n1903_));
  INV_X1    g1461(.A(new_n1898_), .ZN(new_n1904_));
  OAI211_X1 g1462(.A(new_n1176_), .B(new_n1571_), .C1(new_n1904_), .C2(new_n1895_), .ZN(new_n1905_));
  NAND3_X1  g1463(.A1(new_n1905_), .A2(new_n1891_), .A3(new_n1900_), .ZN(new_n1906_));
  NAND3_X1  g1464(.A1(new_n1903_), .A2(new_n1540_), .A3(new_n1906_), .ZN(new_n1907_));
  OAI21_X1  g1465(.A(new_n1891_), .B1(new_n1901_), .B2(new_n1902_), .ZN(new_n1908_));
  NAND4_X1  g1466(.A1(new_n1892_), .A2(new_n1905_), .A3(new_n1900_), .A4(new_n1894_), .ZN(new_n1909_));
  NAND3_X1  g1467(.A1(new_n1908_), .A2(new_n1909_), .A3(new_n680_), .ZN(new_n1910_));
  NAND3_X1  g1468(.A1(new_n1907_), .A2(new_n1910_), .A3(new_n561_), .ZN(new_n1911_));
  NAND2_X1  g1469(.A1(new_n1911_), .A2(new_n577_), .ZN(new_n1912_));
  NAND2_X1  g1470(.A1(new_n1903_), .A2(new_n1906_), .ZN(new_n1913_));
  NAND2_X1  g1471(.A1(new_n1913_), .A2(new_n680_), .ZN(new_n1914_));
  AOI21_X1  g1472(.A(new_n561_), .B1(new_n1914_), .B2(new_n1907_), .ZN(new_n1915_));
  OAI21_X1  g1473(.A(KEYINPUT116), .B1(new_n1912_), .B2(new_n1915_), .ZN(new_n1916_));
  INV_X1    g1474(.A(new_n544_), .ZN(new_n1917_));
  AND3_X1   g1475(.A1(new_n1903_), .A2(new_n1540_), .A3(new_n1906_), .ZN(new_n1918_));
  AOI21_X1  g1476(.A(new_n1540_), .B1(new_n1903_), .B2(new_n1906_), .ZN(new_n1919_));
  INV_X1    g1477(.A(new_n561_), .ZN(new_n1920_));
  NOR3_X1   g1478(.A1(new_n1918_), .A2(new_n1919_), .A3(new_n1920_), .ZN(new_n1921_));
  AOI21_X1  g1479(.A(new_n561_), .B1(new_n1907_), .B2(new_n1910_), .ZN(new_n1922_));
  OAI21_X1  g1480(.A(new_n1917_), .B1(new_n1921_), .B2(new_n1922_), .ZN(new_n1923_));
  OAI21_X1  g1481(.A(new_n1920_), .B1(new_n1918_), .B2(new_n1919_), .ZN(new_n1924_));
  INV_X1    g1482(.A(KEYINPUT116), .ZN(new_n1925_));
  NAND4_X1  g1483(.A1(new_n1924_), .A2(new_n1925_), .A3(new_n577_), .A4(new_n1911_), .ZN(new_n1926_));
  NAND3_X1  g1484(.A1(new_n1916_), .A2(new_n1923_), .A3(new_n1926_), .ZN(new_n1927_));
  NAND2_X1  g1485(.A1(new_n1927_), .A2(new_n564_), .ZN(new_n1928_));
  INV_X1    g1486(.A(new_n1922_), .ZN(new_n1929_));
  NAND3_X1  g1487(.A1(new_n1914_), .A2(new_n561_), .A3(new_n1907_), .ZN(new_n1930_));
  NAND3_X1  g1488(.A1(new_n1929_), .A2(new_n1930_), .A3(new_n544_), .ZN(new_n1931_));
  NAND3_X1  g1489(.A1(new_n1923_), .A2(new_n1182_), .A3(new_n1931_), .ZN(new_n1932_));
  AOI21_X1  g1490(.A(new_n569_), .B1(new_n1928_), .B2(new_n1932_), .ZN(new_n1933_));
  NOR3_X1   g1491(.A1(new_n1921_), .A2(new_n1917_), .A3(new_n1922_), .ZN(new_n1934_));
  AOI21_X1  g1492(.A(new_n544_), .B1(new_n1929_), .B2(new_n1930_), .ZN(new_n1935_));
  OAI21_X1  g1493(.A(new_n1573_), .B1(new_n1934_), .B2(new_n1935_), .ZN(new_n1936_));
  NAND4_X1  g1494(.A1(new_n1916_), .A2(new_n1923_), .A3(new_n563_), .A4(new_n1926_), .ZN(new_n1937_));
  AND3_X1   g1495(.A1(new_n1936_), .A2(new_n1937_), .A3(new_n569_), .ZN(new_n1938_));
  OAI21_X1  g1496(.A(new_n1890_), .B1(new_n1933_), .B2(new_n1938_), .ZN(new_n1939_));
  NAND2_X1  g1497(.A1(new_n529_), .A2(new_n515_), .ZN(new_n1940_));
  INV_X1    g1498(.A(new_n522_), .ZN(new_n1941_));
  OAI21_X1  g1499(.A(new_n1940_), .B1(new_n1941_), .B2(new_n529_), .ZN(new_n1942_));
  XNOR2_X1  g1500(.A(new_n1942_), .B(new_n587_), .ZN(new_n1943_));
  XNOR2_X1  g1501(.A(new_n1943_), .B(new_n586_), .ZN(new_n1944_));
  XNOR2_X1  g1502(.A(new_n1944_), .B(new_n530_), .ZN(new_n1945_));
  NAND2_X1  g1503(.A1(new_n1945_), .A2(new_n1593_), .ZN(new_n1946_));
  OAI21_X1  g1504(.A(new_n1946_), .B1(new_n1587_), .B2(new_n1945_), .ZN(new_n1947_));
  AND2_X1   g1505(.A1(new_n1947_), .A2(new_n520_), .ZN(new_n1948_));
  NOR2_X1   g1506(.A1(new_n1947_), .A2(new_n520_), .ZN(new_n1949_));
  NOR2_X1   g1507(.A1(new_n1948_), .A2(new_n1949_), .ZN(new_n1950_));
  XNOR2_X1  g1508(.A(new_n582_), .B(KEYINPUT117), .ZN(new_n1951_));
  INV_X1    g1509(.A(new_n1184_), .ZN(new_n1952_));
  OAI211_X1 g1510(.A(new_n1950_), .B(new_n1951_), .C1(new_n1952_), .C2(new_n1889_), .ZN(new_n1953_));
  AOI22_X1  g1511(.A1(new_n1591_), .A2(new_n515_), .B1(new_n522_), .B2(new_n1578_), .ZN(new_n1954_));
  XNOR2_X1  g1512(.A(new_n1954_), .B(new_n586_), .ZN(new_n1955_));
  XNOR2_X1  g1513(.A(new_n1955_), .B(new_n587_), .ZN(new_n1956_));
  XNOR2_X1  g1514(.A(new_n1581_), .B(new_n1956_), .ZN(new_n1957_));
  NAND2_X1  g1515(.A1(new_n1957_), .A2(new_n589_), .ZN(new_n1958_));
  OAI21_X1  g1516(.A(new_n1958_), .B1(new_n523_), .B2(new_n1957_), .ZN(new_n1959_));
  XNOR2_X1  g1517(.A(new_n1959_), .B(new_n584_), .ZN(new_n1960_));
  AOI21_X1  g1518(.A(new_n1889_), .B1(new_n1952_), .B2(new_n1951_), .ZN(new_n1961_));
  NOR2_X1   g1519(.A1(new_n1890_), .A2(new_n582_), .ZN(new_n1962_));
  OAI21_X1  g1520(.A(new_n1960_), .B1(new_n1961_), .B2(new_n1962_), .ZN(new_n1963_));
  AND2_X1   g1521(.A1(new_n1953_), .A2(new_n1963_), .ZN(new_n1964_));
  NAND2_X1  g1522(.A1(new_n1555_), .A2(new_n1570_), .ZN(new_n1965_));
  NAND2_X1  g1523(.A1(new_n1554_), .A2(new_n1571_), .ZN(new_n1966_));
  NAND2_X1  g1524(.A1(new_n1965_), .A2(new_n1966_), .ZN(new_n1967_));
  NAND2_X1  g1525(.A1(new_n1967_), .A2(new_n1920_), .ZN(new_n1968_));
  NAND3_X1  g1526(.A1(new_n1965_), .A2(new_n561_), .A3(new_n1966_), .ZN(new_n1969_));
  NOR2_X1   g1527(.A1(new_n553_), .A2(G4394), .ZN(new_n1970_));
  NAND2_X1  g1528(.A1(new_n1560_), .A2(new_n1562_), .ZN(new_n1971_));
  AOI21_X1  g1529(.A(new_n1970_), .B1(new_n1896_), .B2(new_n1971_), .ZN(new_n1972_));
  NAND2_X1  g1530(.A1(new_n1570_), .A2(new_n1182_), .ZN(new_n1973_));
  AOI21_X1  g1531(.A(new_n554_), .B1(new_n1973_), .B2(new_n549_), .ZN(new_n1974_));
  NOR2_X1   g1532(.A1(new_n1972_), .A2(new_n1974_), .ZN(new_n1975_));
  INV_X1    g1533(.A(new_n1975_), .ZN(new_n1976_));
  NAND3_X1  g1534(.A1(new_n1968_), .A2(new_n1969_), .A3(new_n1976_), .ZN(new_n1977_));
  INV_X1    g1535(.A(new_n1977_), .ZN(new_n1978_));
  AOI21_X1  g1536(.A(new_n1976_), .B1(new_n1968_), .B2(new_n1969_), .ZN(new_n1979_));
  NOR3_X1   g1537(.A1(new_n1978_), .A2(new_n1979_), .A3(new_n1917_), .ZN(new_n1980_));
  NAND2_X1  g1538(.A1(new_n1968_), .A2(new_n1969_), .ZN(new_n1981_));
  NAND2_X1  g1539(.A1(new_n1981_), .A2(new_n1975_), .ZN(new_n1982_));
  AOI21_X1  g1540(.A(new_n544_), .B1(new_n1982_), .B2(new_n1977_), .ZN(new_n1983_));
  OAI21_X1  g1541(.A(new_n1573_), .B1(new_n1980_), .B2(new_n1983_), .ZN(new_n1984_));
  NAND3_X1  g1542(.A1(new_n1982_), .A2(new_n1977_), .A3(new_n577_), .ZN(new_n1985_));
  INV_X1    g1543(.A(new_n1985_), .ZN(new_n1986_));
  OAI21_X1  g1544(.A(new_n1917_), .B1(new_n1978_), .B2(new_n1979_), .ZN(new_n1987_));
  NAND2_X1  g1545(.A1(new_n1987_), .A2(new_n563_), .ZN(new_n1988_));
  OAI21_X1  g1546(.A(new_n1984_), .B1(new_n1986_), .B2(new_n1988_), .ZN(new_n1989_));
  INV_X1    g1547(.A(new_n569_), .ZN(new_n1990_));
  AOI21_X1  g1548(.A(new_n1890_), .B1(new_n1989_), .B2(new_n1990_), .ZN(new_n1991_));
  OAI211_X1 g1549(.A(new_n1984_), .B(new_n569_), .C1(new_n1986_), .C2(new_n1988_), .ZN(new_n1992_));
  AOI21_X1  g1550(.A(new_n1964_), .B1(new_n1991_), .B2(new_n1992_), .ZN(new_n1993_));
  INV_X1    g1551(.A(KEYINPUT118), .ZN(new_n1994_));
  AND3_X1   g1552(.A1(new_n1939_), .A2(new_n1993_), .A3(new_n1994_), .ZN(new_n1995_));
  AOI21_X1  g1553(.A(new_n1994_), .B1(new_n1939_), .B2(new_n1993_), .ZN(new_n1996_));
  INV_X1    g1554(.A(new_n1964_), .ZN(new_n1997_));
  AOI21_X1  g1555(.A(new_n569_), .B1(new_n1936_), .B2(new_n1937_), .ZN(new_n1998_));
  OAI21_X1  g1556(.A(new_n1890_), .B1(new_n1938_), .B2(new_n1998_), .ZN(new_n1999_));
  NAND2_X1  g1557(.A1(new_n1991_), .A2(new_n1992_), .ZN(new_n2000_));
  AOI21_X1  g1558(.A(new_n1997_), .B1(new_n1999_), .B2(new_n2000_), .ZN(new_n2001_));
  NOR3_X1   g1559(.A1(new_n1995_), .A2(new_n1996_), .A3(new_n2001_), .ZN(G370));
  NAND2_X1  g1560(.A1(new_n652_), .A2(new_n657_), .ZN(new_n2003_));
  NOR2_X1   g1561(.A1(new_n2003_), .A2(new_n1171_), .ZN(new_n2004_));
  NAND2_X1  g1562(.A1(new_n663_), .A2(new_n2004_), .ZN(new_n2005_));
  INV_X1    g1563(.A(new_n2004_), .ZN(new_n2006_));
  NAND4_X1  g1564(.A1(new_n661_), .A2(new_n2006_), .A3(new_n662_), .A4(new_n1172_), .ZN(new_n2007_));
  OAI21_X1  g1565(.A(new_n503_), .B1(new_n1217_), .B2(new_n1218_), .ZN(new_n2008_));
  NAND2_X1  g1566(.A1(new_n1219_), .A2(new_n1221_), .ZN(new_n2009_));
  OAI21_X1  g1567(.A(new_n2008_), .B1(new_n2009_), .B2(new_n503_), .ZN(new_n2010_));
  AND3_X1   g1568(.A1(new_n2005_), .A2(new_n2007_), .A3(new_n2010_), .ZN(new_n2011_));
  AOI21_X1  g1569(.A(new_n2010_), .B1(new_n2005_), .B2(new_n2007_), .ZN(new_n2012_));
  OAI21_X1  g1570(.A(new_n504_), .B1(new_n2011_), .B2(new_n2012_), .ZN(new_n2013_));
  NAND2_X1  g1571(.A1(new_n2005_), .A2(new_n2007_), .ZN(new_n2014_));
  INV_X1    g1572(.A(new_n2010_), .ZN(new_n2015_));
  NAND2_X1  g1573(.A1(new_n2014_), .A2(new_n2015_), .ZN(new_n2016_));
  NAND3_X1  g1574(.A1(new_n2005_), .A2(new_n2010_), .A3(new_n2007_), .ZN(new_n2017_));
  NAND3_X1  g1575(.A1(new_n2016_), .A2(new_n1202_), .A3(new_n2017_), .ZN(new_n2018_));
  NAND3_X1  g1576(.A1(new_n2013_), .A2(new_n2018_), .A3(KEYINPUT119), .ZN(new_n2019_));
  INV_X1    g1577(.A(KEYINPUT119), .ZN(new_n2020_));
  NAND4_X1  g1578(.A1(new_n2016_), .A2(new_n2020_), .A3(new_n2017_), .A4(new_n1202_), .ZN(new_n2021_));
  NAND3_X1  g1579(.A1(new_n2019_), .A2(new_n1204_), .A3(new_n2021_), .ZN(new_n2022_));
  NAND3_X1  g1580(.A1(new_n2013_), .A2(new_n2018_), .A3(new_n1220_), .ZN(new_n2023_));
  AND3_X1   g1581(.A1(new_n2022_), .A2(new_n670_), .A3(new_n2023_), .ZN(new_n2024_));
  AOI21_X1  g1582(.A(new_n670_), .B1(new_n2022_), .B2(new_n2023_), .ZN(new_n2025_));
  OAI21_X1  g1583(.A(new_n1212_), .B1(new_n2024_), .B2(new_n2025_), .ZN(new_n2026_));
  NAND3_X1  g1584(.A1(new_n2022_), .A2(new_n670_), .A3(new_n2023_), .ZN(new_n2027_));
  NAND3_X1  g1585(.A1(new_n2019_), .A2(new_n1220_), .A3(new_n2021_), .ZN(new_n2028_));
  NAND3_X1  g1586(.A1(new_n2013_), .A2(new_n2018_), .A3(new_n1204_), .ZN(new_n2029_));
  NAND3_X1  g1587(.A1(new_n2028_), .A2(new_n1173_), .A3(new_n2029_), .ZN(new_n2030_));
  NAND3_X1  g1588(.A1(new_n2027_), .A2(new_n2030_), .A3(new_n668_), .ZN(new_n2031_));
  AND3_X1   g1589(.A1(new_n2026_), .A2(new_n635_), .A3(new_n2031_), .ZN(new_n2032_));
  AOI21_X1  g1590(.A(new_n635_), .B1(new_n2026_), .B2(new_n2031_), .ZN(new_n2033_));
  OAI21_X1  g1591(.A(G4526), .B1(new_n2032_), .B2(new_n2033_), .ZN(new_n2034_));
  NAND2_X1  g1592(.A1(new_n2034_), .A2(KEYINPUT127), .ZN(new_n2035_));
  INV_X1    g1593(.A(KEYINPUT127), .ZN(new_n2036_));
  OAI211_X1 g1594(.A(new_n2036_), .B(G4526), .C1(new_n2032_), .C2(new_n2033_), .ZN(new_n2037_));
  INV_X1    g1595(.A(new_n1212_), .ZN(new_n2038_));
  OAI21_X1  g1596(.A(new_n501_), .B1(new_n1217_), .B2(new_n1218_), .ZN(new_n2039_));
  NAND4_X1  g1597(.A1(new_n1231_), .A2(new_n501_), .A3(new_n2038_), .A4(new_n1232_), .ZN(new_n2040_));
  INV_X1    g1598(.A(new_n501_), .ZN(new_n2041_));
  XNOR2_X1  g1599(.A(new_n659_), .B(KEYINPUT59), .ZN(new_n2042_));
  OAI211_X1 g1600(.A(new_n2041_), .B(new_n2042_), .C1(new_n652_), .C2(new_n1212_), .ZN(new_n2043_));
  NAND3_X1  g1601(.A1(new_n2039_), .A2(new_n2040_), .A3(new_n2043_), .ZN(new_n2044_));
  NAND2_X1  g1602(.A1(new_n2044_), .A2(new_n2003_), .ZN(new_n2045_));
  INV_X1    g1603(.A(new_n2003_), .ZN(new_n2046_));
  NAND4_X1  g1604(.A1(new_n2039_), .A2(new_n2040_), .A3(new_n2046_), .A4(new_n2043_), .ZN(new_n2047_));
  AND2_X1   g1605(.A1(new_n2045_), .A2(new_n2047_), .ZN(new_n2048_));
  NAND2_X1  g1606(.A1(new_n663_), .A2(KEYINPUT121), .ZN(new_n2049_));
  INV_X1    g1607(.A(KEYINPUT121), .ZN(new_n2050_));
  NAND3_X1  g1608(.A1(new_n661_), .A2(new_n2050_), .A3(new_n662_), .ZN(new_n2051_));
  NAND4_X1  g1609(.A1(new_n2048_), .A2(KEYINPUT122), .A3(new_n2049_), .A4(new_n2051_), .ZN(new_n2052_));
  INV_X1    g1610(.A(KEYINPUT122), .ZN(new_n2053_));
  NAND2_X1  g1611(.A1(new_n2049_), .A2(new_n2051_), .ZN(new_n2054_));
  NAND2_X1  g1612(.A1(new_n2045_), .A2(new_n2047_), .ZN(new_n2055_));
  OAI21_X1  g1613(.A(new_n2053_), .B1(new_n2054_), .B2(new_n2055_), .ZN(new_n2056_));
  NAND2_X1  g1614(.A1(new_n2052_), .A2(new_n2056_), .ZN(new_n2057_));
  NAND2_X1  g1615(.A1(new_n2055_), .A2(new_n663_), .ZN(new_n2058_));
  INV_X1    g1616(.A(KEYINPUT120), .ZN(new_n2059_));
  NAND2_X1  g1617(.A1(new_n2058_), .A2(new_n2059_), .ZN(new_n2060_));
  NAND3_X1  g1618(.A1(new_n2055_), .A2(KEYINPUT120), .A3(new_n663_), .ZN(new_n2061_));
  NAND2_X1  g1619(.A1(new_n2060_), .A2(new_n2061_), .ZN(new_n2062_));
  NAND2_X1  g1620(.A1(new_n2057_), .A2(new_n2062_), .ZN(new_n2063_));
  NAND2_X1  g1621(.A1(new_n2063_), .A2(new_n1202_), .ZN(new_n2064_));
  NAND3_X1  g1622(.A1(new_n2057_), .A2(new_n2062_), .A3(new_n504_), .ZN(new_n2065_));
  AOI21_X1  g1623(.A(new_n1220_), .B1(new_n2064_), .B2(new_n2065_), .ZN(new_n2066_));
  AOI22_X1  g1624(.A1(new_n2049_), .A2(new_n2051_), .B1(new_n2045_), .B2(new_n2047_), .ZN(new_n2067_));
  INV_X1    g1625(.A(KEYINPUT123), .ZN(new_n2068_));
  OAI22_X1  g1626(.A1(new_n2067_), .A2(new_n2068_), .B1(new_n663_), .B2(new_n2055_), .ZN(new_n2069_));
  AND2_X1   g1627(.A1(new_n2067_), .A2(new_n2068_), .ZN(new_n2070_));
  OAI21_X1  g1628(.A(new_n1202_), .B1(new_n2069_), .B2(new_n2070_), .ZN(new_n2071_));
  AND3_X1   g1629(.A1(new_n2065_), .A2(new_n2071_), .A3(new_n1220_), .ZN(new_n2072_));
  OAI21_X1  g1630(.A(new_n1173_), .B1(new_n2066_), .B2(new_n2072_), .ZN(new_n2073_));
  AND3_X1   g1631(.A1(new_n2057_), .A2(new_n2062_), .A3(new_n504_), .ZN(new_n2074_));
  AOI21_X1  g1632(.A(new_n504_), .B1(new_n2057_), .B2(new_n2062_), .ZN(new_n2075_));
  OAI21_X1  g1633(.A(new_n1204_), .B1(new_n2074_), .B2(new_n2075_), .ZN(new_n2076_));
  NAND3_X1  g1634(.A1(new_n2065_), .A2(new_n2071_), .A3(new_n1220_), .ZN(new_n2077_));
  NAND3_X1  g1635(.A1(new_n2076_), .A2(new_n670_), .A3(new_n2077_), .ZN(new_n2078_));
  AOI21_X1  g1636(.A(new_n2038_), .B1(new_n2073_), .B2(new_n2078_), .ZN(new_n2079_));
  INV_X1    g1637(.A(KEYINPUT124), .ZN(new_n2080_));
  NAND3_X1  g1638(.A1(new_n2065_), .A2(new_n2071_), .A3(new_n1204_), .ZN(new_n2081_));
  NAND2_X1  g1639(.A1(new_n2081_), .A2(new_n1173_), .ZN(new_n2082_));
  AOI21_X1  g1640(.A(new_n1204_), .B1(new_n2064_), .B2(new_n2065_), .ZN(new_n2083_));
  OAI21_X1  g1641(.A(new_n668_), .B1(new_n2082_), .B2(new_n2083_), .ZN(new_n2084_));
  AND3_X1   g1642(.A1(new_n2076_), .A2(new_n670_), .A3(new_n2077_), .ZN(new_n2085_));
  OAI21_X1  g1643(.A(new_n2080_), .B1(new_n2084_), .B2(new_n2085_), .ZN(new_n2086_));
  OAI21_X1  g1644(.A(new_n1220_), .B1(new_n2074_), .B2(new_n2075_), .ZN(new_n2087_));
  NAND3_X1  g1645(.A1(new_n2087_), .A2(new_n1173_), .A3(new_n2081_), .ZN(new_n2088_));
  NAND4_X1  g1646(.A1(new_n2078_), .A2(new_n2088_), .A3(KEYINPUT124), .A4(new_n668_), .ZN(new_n2089_));
  AOI21_X1  g1647(.A(new_n2079_), .B1(new_n2086_), .B2(new_n2089_), .ZN(new_n2090_));
  OAI21_X1  g1648(.A(new_n505_), .B1(new_n2090_), .B2(new_n635_), .ZN(new_n2091_));
  AOI211_X1 g1649(.A(new_n1203_), .B(new_n2079_), .C1(new_n2086_), .C2(new_n2089_), .ZN(new_n2092_));
  OAI211_X1 g1650(.A(new_n2035_), .B(new_n2037_), .C1(new_n2091_), .C2(new_n2092_), .ZN(new_n2093_));
  NOR2_X1   g1651(.A1(new_n607_), .A2(new_n674_), .ZN(new_n2094_));
  INV_X1    g1652(.A(new_n2094_), .ZN(new_n2095_));
  AOI21_X1  g1653(.A(new_n610_), .B1(new_n1238_), .B2(new_n2095_), .ZN(new_n2096_));
  XNOR2_X1  g1654(.A(new_n1241_), .B(new_n2096_), .ZN(new_n2097_));
  XNOR2_X1  g1655(.A(new_n673_), .B(new_n675_), .ZN(new_n2098_));
  XNOR2_X1  g1656(.A(new_n2097_), .B(new_n2098_), .ZN(new_n2099_));
  NOR2_X1   g1657(.A1(new_n2099_), .A2(new_n603_), .ZN(new_n2100_));
  NAND2_X1  g1658(.A1(new_n2099_), .A2(new_n603_), .ZN(new_n2101_));
  AOI21_X1  g1659(.A(new_n2100_), .B1(KEYINPUT125), .B2(new_n2101_), .ZN(new_n2102_));
  OAI21_X1  g1660(.A(new_n2102_), .B1(KEYINPUT125), .B2(new_n2101_), .ZN(new_n2103_));
  NOR2_X1   g1661(.A1(new_n665_), .A2(G4526), .ZN(new_n2104_));
  INV_X1    g1662(.A(new_n1888_), .ZN(new_n2105_));
  AND2_X1   g1663(.A1(new_n607_), .A2(new_n674_), .ZN(new_n2106_));
  OAI21_X1  g1664(.A(new_n614_), .B1(new_n2106_), .B2(new_n2094_), .ZN(new_n2107_));
  NAND2_X1  g1665(.A1(new_n2107_), .A2(new_n1250_), .ZN(new_n2108_));
  XNOR2_X1  g1666(.A(new_n2108_), .B(new_n673_), .ZN(new_n2109_));
  XNOR2_X1  g1667(.A(new_n2109_), .B(new_n610_), .ZN(new_n2110_));
  INV_X1    g1668(.A(new_n603_), .ZN(new_n2111_));
  NOR3_X1   g1669(.A1(new_n1251_), .A2(new_n617_), .A3(new_n2111_), .ZN(new_n2112_));
  AOI21_X1  g1670(.A(new_n2112_), .B1(new_n2111_), .B2(new_n617_), .ZN(new_n2113_));
  XNOR2_X1  g1671(.A(new_n2110_), .B(new_n2113_), .ZN(new_n2114_));
  AOI22_X1  g1672(.A1(new_n2103_), .A2(new_n2104_), .B1(new_n2105_), .B2(new_n2114_), .ZN(new_n2115_));
  NAND3_X1  g1673(.A1(new_n665_), .A2(KEYINPUT126), .A3(new_n1887_), .ZN(new_n2116_));
  INV_X1    g1674(.A(KEYINPUT126), .ZN(new_n2117_));
  INV_X1    g1675(.A(new_n665_), .ZN(new_n2118_));
  OAI21_X1  g1676(.A(new_n2117_), .B1(new_n2118_), .B2(new_n1174_), .ZN(new_n2119_));
  NAND4_X1  g1677(.A1(new_n2103_), .A2(G4526), .A3(new_n2116_), .A4(new_n2119_), .ZN(new_n2120_));
  AND2_X1   g1678(.A1(new_n2115_), .A2(new_n2120_), .ZN(new_n2121_));
  AND2_X1   g1679(.A1(new_n2086_), .A2(new_n2089_), .ZN(new_n2122_));
  OAI21_X1  g1680(.A(new_n1203_), .B1(new_n2122_), .B2(new_n2079_), .ZN(new_n2123_));
  NAND2_X1  g1681(.A1(new_n2090_), .A2(new_n635_), .ZN(new_n2124_));
  NAND3_X1  g1682(.A1(new_n2123_), .A2(new_n505_), .A3(new_n2124_), .ZN(new_n2125_));
  INV_X1    g1683(.A(new_n2032_), .ZN(new_n2126_));
  NOR3_X1   g1684(.A1(new_n2024_), .A2(new_n2025_), .A3(new_n1212_), .ZN(new_n2127_));
  AOI21_X1  g1685(.A(new_n668_), .B1(new_n2030_), .B2(new_n2027_), .ZN(new_n2128_));
  OAI21_X1  g1686(.A(new_n1203_), .B1(new_n2127_), .B2(new_n2128_), .ZN(new_n2129_));
  NAND2_X1  g1687(.A1(new_n2126_), .A2(new_n2129_), .ZN(new_n2130_));
  AOI21_X1  g1688(.A(new_n2121_), .B1(new_n2130_), .B2(G4526), .ZN(new_n2131_));
  AOI22_X1  g1689(.A1(new_n2093_), .A2(new_n2121_), .B1(new_n2125_), .B2(new_n2131_), .ZN(G399));
endmodule


