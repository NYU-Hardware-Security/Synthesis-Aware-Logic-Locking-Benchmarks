//Secret key is'0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_c1355" written by ABC on Wed Oct 26 13:34:58 2022

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n470_, new_n471_, new_n472_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n520_, new_n521_,
    new_n522_, new_n524_, new_n525_, new_n526_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n626_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n640_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n138_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n139_));
  NAND2_X1  g002(.A1(new_n139_), .A2(KEYINPUT25), .ZN(new_n140_));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n141_));
  NAND3_X1  g004(.A1(new_n141_), .A2(G183gat), .A3(G190gat), .ZN(new_n142_));
  INV_X1    g005(.A(G183gat), .ZN(new_n143_));
  INV_X1    g006(.A(G190gat), .ZN(new_n144_));
  NAND2_X1  g007(.A1(new_n143_), .A2(new_n144_), .ZN(new_n145_));
  NAND3_X1  g008(.A1(new_n140_), .A2(new_n142_), .A3(new_n145_), .ZN(new_n146_));
  INV_X1    g009(.A(G169gat), .ZN(new_n147_));
  INV_X1    g010(.A(G176gat), .ZN(new_n148_));
  NAND3_X1  g011(.A1(new_n147_), .A2(new_n148_), .A3(KEYINPUT24), .ZN(new_n149_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n150_));
  OAI21_X1  g013(.A(new_n150_), .B1(G169gat), .B2(G176gat), .ZN(new_n151_));
  NAND2_X1  g014(.A1(new_n149_), .A2(new_n151_), .ZN(new_n152_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n153_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n154_));
  NAND2_X1  g017(.A1(new_n153_), .A2(new_n154_), .ZN(new_n155_));
  NAND3_X1  g018(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n156_));
  NAND2_X1  g019(.A1(new_n155_), .A2(new_n156_), .ZN(new_n157_));
  NAND3_X1  g020(.A1(new_n146_), .A2(new_n152_), .A3(new_n157_), .ZN(new_n158_));
  NAND2_X1  g021(.A1(new_n144_), .A2(KEYINPUT26), .ZN(new_n159_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n160_));
  NAND2_X1  g023(.A1(new_n160_), .A2(G190gat), .ZN(new_n161_));
  NAND3_X1  g024(.A1(new_n159_), .A2(new_n161_), .A3(new_n143_), .ZN(new_n162_));
  XNOR2_X1  g025(.A(G169gat), .B(G176gat), .ZN(new_n163_));
  NAND3_X1  g026(.A1(new_n162_), .A2(new_n139_), .A3(new_n163_), .ZN(new_n164_));
  NAND2_X1  g027(.A1(new_n158_), .A2(new_n164_), .ZN(new_n165_));
  INV_X1    g028(.A(G134gat), .ZN(new_n166_));
  NAND2_X1  g029(.A1(new_n166_), .A2(G127gat), .ZN(new_n167_));
  INV_X1    g030(.A(G127gat), .ZN(new_n168_));
  NAND2_X1  g031(.A1(new_n168_), .A2(G134gat), .ZN(new_n169_));
  NAND2_X1  g032(.A1(new_n167_), .A2(new_n169_), .ZN(new_n170_));
  INV_X1    g033(.A(G120gat), .ZN(new_n171_));
  NAND2_X1  g034(.A1(new_n171_), .A2(G113gat), .ZN(new_n172_));
  INV_X1    g035(.A(G113gat), .ZN(new_n173_));
  NAND2_X1  g036(.A1(new_n173_), .A2(G120gat), .ZN(new_n174_));
  NAND2_X1  g037(.A1(new_n172_), .A2(new_n174_), .ZN(new_n175_));
  NAND3_X1  g038(.A1(new_n170_), .A2(new_n175_), .A3(KEYINPUT1), .ZN(new_n176_));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n177_));
  NAND3_X1  g040(.A1(new_n167_), .A2(new_n169_), .A3(new_n177_), .ZN(new_n178_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n179_));
  NAND2_X1  g042(.A1(new_n178_), .A2(new_n179_), .ZN(new_n180_));
  AOI21_X1  g043(.A(new_n177_), .B1(new_n167_), .B2(new_n169_), .ZN(new_n181_));
  OAI21_X1  g044(.A(new_n176_), .B1(new_n180_), .B2(new_n181_), .ZN(new_n182_));
  NAND2_X1  g045(.A1(new_n182_), .A2(KEYINPUT4), .ZN(new_n183_));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n184_));
  OAI211_X1 g047(.A(new_n176_), .B(new_n184_), .C1(new_n180_), .C2(new_n181_), .ZN(new_n185_));
  INV_X1    g048(.A(G227gat), .ZN(new_n186_));
  INV_X1    g049(.A(G233gat), .ZN(new_n187_));
  NOR2_X1   g050(.A1(new_n186_), .A2(new_n187_), .ZN(new_n188_));
  INV_X1    g051(.A(new_n188_), .ZN(new_n189_));
  NAND3_X1  g052(.A1(new_n183_), .A2(new_n185_), .A3(new_n189_), .ZN(new_n190_));
  INV_X1    g053(.A(new_n190_), .ZN(new_n191_));
  AOI21_X1  g054(.A(new_n189_), .B1(new_n183_), .B2(new_n185_), .ZN(new_n192_));
  OAI21_X1  g055(.A(new_n165_), .B1(new_n191_), .B2(new_n192_), .ZN(new_n193_));
  INV_X1    g056(.A(new_n192_), .ZN(new_n194_));
  INV_X1    g057(.A(new_n165_), .ZN(new_n195_));
  NAND3_X1  g058(.A1(new_n194_), .A2(new_n195_), .A3(new_n190_), .ZN(new_n196_));
  INV_X1    g059(.A(KEYINPUT31), .ZN(new_n197_));
  NAND3_X1  g060(.A1(new_n193_), .A2(new_n196_), .A3(new_n197_), .ZN(new_n198_));
  XOR2_X1   g061(.A(G15gat), .B(G43gat), .Z(new_n199_));
  NAND2_X1  g062(.A1(new_n198_), .A2(new_n199_), .ZN(new_n200_));
  INV_X1    g063(.A(new_n199_), .ZN(new_n201_));
  NAND4_X1  g064(.A1(new_n193_), .A2(new_n196_), .A3(new_n197_), .A4(new_n201_), .ZN(new_n202_));
  AOI21_X1  g065(.A(new_n138_), .B1(new_n200_), .B2(new_n202_), .ZN(new_n203_));
  INV_X1    g066(.A(new_n203_), .ZN(new_n204_));
  NAND3_X1  g067(.A1(new_n200_), .A2(new_n202_), .A3(new_n138_), .ZN(new_n205_));
  NAND2_X1  g068(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n207_));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n208_));
  XOR2_X1   g071(.A(new_n207_), .B(new_n208_), .Z(new_n209_));
  INV_X1    g072(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g073(.A(G148gat), .ZN(new_n211_));
  NAND2_X1  g074(.A1(new_n211_), .A2(G141gat), .ZN(new_n212_));
  INV_X1    g075(.A(G141gat), .ZN(new_n213_));
  NAND2_X1  g076(.A1(new_n213_), .A2(G148gat), .ZN(new_n214_));
  NAND2_X1  g077(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g078(.A(G155gat), .ZN(new_n216_));
  INV_X1    g079(.A(G162gat), .ZN(new_n217_));
  NAND2_X1  g080(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g081(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NAND2_X1  g082(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g083(.A(KEYINPUT3), .B1(new_n215_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g084(.A(G141gat), .B(G148gat), .ZN(new_n222_));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n223_));
  NAND4_X1  g086(.A1(new_n222_), .A2(new_n223_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n224_));
  NAND3_X1  g087(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT2), .ZN(new_n225_));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n226_));
  OAI21_X1  g089(.A(new_n226_), .B1(G155gat), .B2(G162gat), .ZN(new_n227_));
  NAND3_X1  g090(.A1(new_n225_), .A2(new_n227_), .A3(new_n219_), .ZN(new_n228_));
  AOI22_X1  g091(.A1(new_n221_), .A2(new_n224_), .B1(new_n215_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g092(.A(new_n229_), .B1(new_n183_), .B2(new_n185_), .ZN(new_n230_));
  NAND2_X1  g093(.A1(new_n221_), .A2(new_n224_), .ZN(new_n231_));
  NAND2_X1  g094(.A1(new_n228_), .A2(new_n215_), .ZN(new_n232_));
  NAND2_X1  g095(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g096(.A(new_n182_), .ZN(new_n234_));
  NOR2_X1   g097(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g099(.A(new_n236_), .ZN(new_n237_));
  NOR3_X1   g100(.A1(new_n230_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g101(.A(new_n236_), .B(KEYINPUT0), .ZN(new_n239_));
  INV_X1    g102(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g103(.A1(new_n233_), .A2(new_n234_), .ZN(new_n241_));
  NAND2_X1  g104(.A1(new_n229_), .A2(new_n182_), .ZN(new_n242_));
  AOI21_X1  g105(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g106(.A(new_n210_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g107(.A1(new_n183_), .A2(new_n185_), .ZN(new_n245_));
  NAND2_X1  g108(.A1(new_n245_), .A2(new_n233_), .ZN(new_n246_));
  NAND3_X1  g109(.A1(new_n246_), .A2(new_n242_), .A3(new_n236_), .ZN(new_n247_));
  NAND2_X1  g110(.A1(new_n241_), .A2(new_n242_), .ZN(new_n248_));
  NAND2_X1  g111(.A1(new_n248_), .A2(new_n239_), .ZN(new_n249_));
  NAND3_X1  g112(.A1(new_n247_), .A2(new_n249_), .A3(new_n209_), .ZN(new_n250_));
  NAND2_X1  g113(.A1(new_n244_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g114(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g115(.A(G211gat), .ZN(new_n253_));
  INV_X1    g116(.A(G218gat), .ZN(new_n254_));
  NAND3_X1  g117(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT21), .ZN(new_n255_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n256_));
  OAI21_X1  g119(.A(new_n256_), .B1(G211gat), .B2(G218gat), .ZN(new_n257_));
  NAND2_X1  g120(.A1(G211gat), .A2(G218gat), .ZN(new_n258_));
  NAND3_X1  g121(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XOR2_X1   g122(.A(G197gat), .B(G204gat), .Z(new_n260_));
  NAND2_X1  g123(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g124(.A1(new_n254_), .A2(KEYINPUT22), .ZN(new_n262_));
  INV_X1    g125(.A(KEYINPUT22), .ZN(new_n263_));
  NAND2_X1  g126(.A1(new_n263_), .A2(G218gat), .ZN(new_n264_));
  NAND3_X1  g127(.A1(new_n262_), .A2(new_n264_), .A3(new_n253_), .ZN(new_n265_));
  XNOR2_X1  g128(.A(G197gat), .B(G204gat), .ZN(new_n266_));
  NAND3_X1  g129(.A1(new_n265_), .A2(new_n266_), .A3(new_n258_), .ZN(new_n267_));
  NAND2_X1  g130(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g131(.A(new_n233_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n270_));
  INV_X1    g133(.A(new_n270_), .ZN(new_n271_));
  OR2_X1    g134(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g135(.A1(new_n269_), .A2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g136(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g137(.A(G78gat), .B(G106gat), .ZN(new_n275_));
  XNOR2_X1  g138(.A(new_n275_), .B(KEYINPUT29), .ZN(new_n276_));
  XOR2_X1   g139(.A(G22gat), .B(G50gat), .Z(new_n277_));
  XNOR2_X1  g140(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NOR2_X1   g141(.A1(new_n269_), .A2(new_n271_), .ZN(new_n279_));
  OAI21_X1  g142(.A(new_n278_), .B1(new_n279_), .B2(KEYINPUT30), .ZN(new_n280_));
  NAND2_X1  g143(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g144(.A1(new_n272_), .A2(KEYINPUT30), .A3(new_n273_), .A4(new_n278_), .ZN(new_n282_));
  NAND2_X1  g145(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n285_));
  XNOR2_X1  g148(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g149(.A(new_n286_), .B(KEYINPUT20), .ZN(new_n287_));
  INV_X1    g150(.A(new_n287_), .ZN(new_n288_));
  AND2_X1   g151(.A1(G226gat), .A2(G233gat), .ZN(new_n289_));
  NAND4_X1  g152(.A1(new_n158_), .A2(new_n261_), .A3(new_n267_), .A4(new_n164_), .ZN(new_n290_));
  AOI21_X1  g153(.A(new_n289_), .B1(new_n290_), .B2(KEYINPUT27), .ZN(new_n291_));
  NAND2_X1  g154(.A1(new_n165_), .A2(new_n268_), .ZN(new_n292_));
  NAND2_X1  g155(.A1(new_n292_), .A2(new_n290_), .ZN(new_n293_));
  NAND2_X1  g156(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g157(.A(new_n292_), .B(new_n290_), .C1(KEYINPUT27), .C2(new_n289_), .ZN(new_n295_));
  AOI21_X1  g158(.A(new_n288_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g159(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g160(.A1(new_n288_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n298_));
  NAND2_X1  g161(.A1(new_n298_), .A2(KEYINPUT28), .ZN(new_n299_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n300_));
  NAND4_X1  g163(.A1(new_n288_), .A2(new_n294_), .A3(new_n300_), .A4(new_n295_), .ZN(new_n301_));
  NAND3_X1  g164(.A1(new_n297_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  NOR2_X1   g165(.A1(new_n283_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g166(.A1(new_n206_), .A2(new_n252_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g167(.A(KEYINPUT35), .ZN(new_n305_));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n306_));
  AND3_X1   g169(.A1(new_n294_), .A2(new_n306_), .A3(new_n295_), .ZN(new_n307_));
  AOI21_X1  g170(.A(new_n306_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n308_));
  OAI21_X1  g171(.A(new_n286_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g172(.A1(new_n309_), .A2(KEYINPUT34), .ZN(new_n310_));
  INV_X1    g173(.A(KEYINPUT34), .ZN(new_n311_));
  OAI211_X1 g174(.A(new_n311_), .B(new_n286_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n312_));
  AOI21_X1  g175(.A(new_n296_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n313_));
  NAND3_X1  g176(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g177(.A(new_n236_), .B1(new_n246_), .B2(new_n242_), .ZN(new_n315_));
  NOR2_X1   g178(.A1(new_n248_), .A2(new_n239_), .ZN(new_n316_));
  OAI21_X1  g179(.A(new_n210_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g180(.A1(new_n302_), .A2(new_n250_), .A3(new_n317_), .ZN(new_n318_));
  AND2_X1   g181(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g182(.A(new_n305_), .B1(new_n319_), .B2(new_n283_), .ZN(new_n320_));
  AOI21_X1  g183(.A(new_n283_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n321_));
  NAND2_X1  g184(.A1(new_n321_), .A2(KEYINPUT35), .ZN(new_n322_));
  INV_X1    g185(.A(new_n302_), .ZN(new_n323_));
  NAND3_X1  g186(.A1(new_n283_), .A2(new_n252_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g187(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g188(.A(KEYINPUT32), .ZN(new_n326_));
  INV_X1    g189(.A(new_n205_), .ZN(new_n327_));
  OAI21_X1  g190(.A(new_n326_), .B1(new_n327_), .B2(new_n203_), .ZN(new_n328_));
  NAND3_X1  g191(.A1(new_n204_), .A2(KEYINPUT32), .A3(new_n205_), .ZN(new_n329_));
  NAND2_X1  g192(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g193(.A(KEYINPUT36), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g194(.A(new_n324_), .B1(new_n321_), .B2(KEYINPUT35), .ZN(new_n332_));
  AOI211_X1 g195(.A(new_n305_), .B(new_n283_), .C1(new_n314_), .C2(new_n318_), .ZN(new_n333_));
  OAI211_X1 g196(.A(new_n330_), .B(KEYINPUT36), .C1(new_n332_), .C2(new_n333_), .ZN(new_n334_));
  INV_X1    g197(.A(new_n334_), .ZN(new_n335_));
  OAI21_X1  g198(.A(new_n304_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g199(.A(G134gat), .B(G162gat), .ZN(new_n337_));
  NAND2_X1  g200(.A1(G232gat), .A2(G233gat), .ZN(new_n338_));
  XOR2_X1   g201(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g202(.A(new_n339_), .ZN(new_n340_));
  XOR2_X1   g203(.A(G99gat), .B(G106gat), .Z(new_n341_));
  INV_X1    g204(.A(G85gat), .ZN(new_n342_));
  INV_X1    g205(.A(G92gat), .ZN(new_n343_));
  NOR2_X1   g206(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g207(.A1(G85gat), .A2(G92gat), .ZN(new_n345_));
  OAI21_X1  g208(.A(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g209(.A(new_n346_), .B(KEYINPUT9), .ZN(new_n347_));
  NAND2_X1  g210(.A1(new_n341_), .A2(KEYINPUT8), .ZN(new_n348_));
  NOR3_X1   g211(.A1(KEYINPUT8), .A2(G99gat), .A3(G106gat), .ZN(new_n349_));
  NOR2_X1   g212(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g213(.A1(new_n345_), .A2(KEYINPUT7), .ZN(new_n351_));
  OR2_X1    g214(.A1(new_n345_), .A2(KEYINPUT7), .ZN(new_n352_));
  NAND4_X1  g215(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g216(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g217(.A(KEYINPUT11), .ZN(new_n355_));
  NAND2_X1  g218(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g219(.A(KEYINPUT15), .ZN(new_n357_));
  AOI21_X1  g220(.A(G36gat), .B1(new_n357_), .B2(G29gat), .ZN(new_n358_));
  OAI21_X1  g221(.A(new_n358_), .B1(new_n357_), .B2(G29gat), .ZN(new_n359_));
  INV_X1    g222(.A(G29gat), .ZN(new_n360_));
  NAND3_X1  g223(.A1(new_n360_), .A2(KEYINPUT15), .A3(G36gat), .ZN(new_n361_));
  NAND2_X1  g224(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g225(.A(G43gat), .B(G50gat), .ZN(new_n363_));
  XNOR2_X1  g226(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND3_X1  g227(.A1(new_n347_), .A2(KEYINPUT11), .A3(new_n353_), .ZN(new_n365_));
  NAND3_X1  g228(.A1(new_n356_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  OR2_X1    g229(.A1(new_n366_), .A2(KEYINPUT37), .ZN(new_n367_));
  XOR2_X1   g230(.A(G190gat), .B(G218gat), .Z(new_n368_));
  INV_X1    g231(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g232(.A1(new_n354_), .A2(new_n364_), .ZN(new_n370_));
  OAI21_X1  g233(.A(new_n366_), .B1(KEYINPUT37), .B2(new_n370_), .ZN(new_n371_));
  AND3_X1   g234(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g235(.A(new_n369_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n373_));
  OAI21_X1  g236(.A(new_n340_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g237(.A1(new_n367_), .A2(new_n371_), .ZN(new_n375_));
  NAND2_X1  g238(.A1(new_n375_), .A2(new_n368_), .ZN(new_n376_));
  NAND3_X1  g239(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n377_));
  NAND3_X1  g240(.A1(new_n376_), .A2(new_n339_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g241(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g242(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g243(.A(G57gat), .B(G64gat), .ZN(new_n381_));
  INV_X1    g244(.A(G78gat), .ZN(new_n382_));
  OR2_X1    g245(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g246(.A(G71gat), .ZN(new_n384_));
  NAND3_X1  g247(.A1(new_n381_), .A2(KEYINPUT10), .A3(new_n382_), .ZN(new_n385_));
  NAND3_X1  g248(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g249(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g250(.A(new_n384_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n388_));
  NOR2_X1   g251(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g252(.A1(new_n389_), .A2(KEYINPUT12), .ZN(new_n390_));
  INV_X1    g253(.A(new_n388_), .ZN(new_n391_));
  NAND2_X1  g254(.A1(new_n391_), .A2(new_n386_), .ZN(new_n392_));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n393_));
  NAND2_X1  g256(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g257(.A1(new_n356_), .A2(new_n390_), .A3(new_n394_), .A4(new_n365_), .ZN(new_n395_));
  NAND2_X1  g258(.A1(G230gat), .A2(G233gat), .ZN(new_n396_));
  OAI21_X1  g259(.A(KEYINPUT13), .B1(new_n354_), .B2(new_n392_), .ZN(new_n397_));
  INV_X1    g260(.A(new_n354_), .ZN(new_n398_));
  INV_X1    g261(.A(KEYINPUT13), .ZN(new_n399_));
  NAND3_X1  g262(.A1(new_n398_), .A2(new_n389_), .A3(new_n399_), .ZN(new_n400_));
  NAND4_X1  g263(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .A4(new_n400_), .ZN(new_n401_));
  INV_X1    g264(.A(new_n396_), .ZN(new_n402_));
  NOR2_X1   g265(.A1(new_n398_), .A2(new_n389_), .ZN(new_n403_));
  NOR2_X1   g266(.A1(new_n354_), .A2(new_n392_), .ZN(new_n404_));
  OAI21_X1  g267(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g268(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g269(.A(G120gat), .B(G148gat), .ZN(new_n407_));
  XNOR2_X1  g270(.A(new_n407_), .B(KEYINPUT5), .ZN(new_n408_));
  XNOR2_X1  g271(.A(G176gat), .B(G204gat), .ZN(new_n409_));
  XNOR2_X1  g272(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XOR2_X1   g273(.A(new_n410_), .B(KEYINPUT6), .Z(new_n411_));
  NAND2_X1  g274(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g275(.A(new_n411_), .ZN(new_n413_));
  NAND3_X1  g276(.A1(new_n401_), .A2(new_n405_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g277(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g278(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n417_));
  INV_X1    g280(.A(new_n364_), .ZN(new_n418_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n419_));
  AND2_X1   g282(.A1(G15gat), .A2(G22gat), .ZN(new_n420_));
  OAI21_X1  g283(.A(new_n419_), .B1(KEYINPUT16), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g284(.A1(G15gat), .A2(G22gat), .ZN(new_n422_));
  NOR2_X1   g285(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g286(.A(new_n421_), .B(new_n423_), .ZN(new_n424_));
  OAI21_X1  g287(.A(new_n417_), .B1(new_n418_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g288(.A(new_n364_), .B(new_n424_), .ZN(new_n426_));
  OAI21_X1  g289(.A(new_n425_), .B1(new_n426_), .B2(new_n417_), .ZN(new_n427_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g291(.A(new_n428_), .B(KEYINPUT14), .ZN(new_n429_));
  NAND2_X1  g292(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g293(.A1(new_n426_), .A2(new_n428_), .ZN(new_n431_));
  NAND2_X1  g294(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g295(.A(G113gat), .B(G141gat), .ZN(new_n433_));
  XNOR2_X1  g296(.A(G169gat), .B(G197gat), .ZN(new_n434_));
  XOR2_X1   g297(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  INV_X1    g298(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g299(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g300(.A1(new_n430_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n438_));
  NAND2_X1  g301(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g302(.A1(new_n416_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g303(.A1(new_n390_), .A2(new_n394_), .ZN(new_n441_));
  OR2_X1    g304(.A1(new_n441_), .A2(new_n424_), .ZN(new_n442_));
  INV_X1    g305(.A(G231gat), .ZN(new_n443_));
  NOR3_X1   g306(.A1(new_n443_), .A2(new_n187_), .A3(KEYINPUT18), .ZN(new_n444_));
  AOI21_X1  g307(.A(new_n444_), .B1(new_n389_), .B2(new_n424_), .ZN(new_n445_));
  XNOR2_X1  g308(.A(G127gat), .B(G155gat), .ZN(new_n446_));
  OAI21_X1  g309(.A(KEYINPUT18), .B1(new_n443_), .B2(new_n187_), .ZN(new_n447_));
  XNOR2_X1  g310(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g311(.A(new_n448_), .ZN(new_n449_));
  AND3_X1   g312(.A1(new_n442_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g313(.A(new_n449_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n451_));
  XNOR2_X1  g314(.A(G183gat), .B(G211gat), .ZN(new_n452_));
  XNOR2_X1  g315(.A(new_n452_), .B(KEYINPUT19), .ZN(new_n453_));
  INV_X1    g316(.A(new_n453_), .ZN(new_n454_));
  OR3_X1    g317(.A1(new_n450_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g318(.A(new_n454_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n456_));
  NAND2_X1  g319(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g320(.A1(new_n440_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g321(.A1(new_n336_), .A2(new_n380_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g322(.A(G1gat), .ZN(new_n460_));
  NOR3_X1   g323(.A1(new_n459_), .A2(new_n460_), .A3(new_n252_), .ZN(new_n461_));
  NOR2_X1   g324(.A1(new_n457_), .A2(new_n379_), .ZN(new_n462_));
  NAND3_X1  g325(.A1(new_n336_), .A2(new_n439_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g326(.A(KEYINPUT38), .ZN(new_n464_));
  NAND2_X1  g327(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g328(.A1(new_n336_), .A2(KEYINPUT38), .A3(new_n439_), .A4(new_n462_), .ZN(new_n466_));
  AND3_X1   g329(.A1(new_n465_), .A2(new_n466_), .A3(new_n416_), .ZN(new_n467_));
  NAND2_X1  g330(.A1(new_n467_), .A2(new_n251_), .ZN(new_n468_));
  AOI21_X1  g331(.A(new_n461_), .B1(new_n468_), .B2(new_n460_), .ZN(G1324gat));
  INV_X1    g332(.A(G8gat), .ZN(new_n470_));
  NOR3_X1   g333(.A1(new_n459_), .A2(new_n470_), .A3(new_n323_), .ZN(new_n471_));
  NAND2_X1  g334(.A1(new_n467_), .A2(new_n302_), .ZN(new_n472_));
  AOI21_X1  g335(.A(new_n471_), .B1(new_n472_), .B2(new_n470_), .ZN(G1325gat));
  INV_X1    g336(.A(new_n206_), .ZN(new_n474_));
  NOR2_X1   g337(.A1(new_n474_), .A2(G15gat), .ZN(new_n475_));
  NAND4_X1  g338(.A1(new_n465_), .A2(new_n466_), .A3(new_n416_), .A4(new_n475_), .ZN(new_n476_));
  OAI21_X1  g339(.A(G15gat), .B1(new_n459_), .B2(new_n330_), .ZN(new_n477_));
  NAND2_X1  g340(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g341(.A(KEYINPUT39), .ZN(new_n479_));
  NAND2_X1  g342(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g343(.A1(new_n476_), .A2(KEYINPUT39), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g344(.A1(new_n480_), .A2(new_n481_), .ZN(G1326gat));
  INV_X1    g345(.A(G22gat), .ZN(new_n483_));
  INV_X1    g346(.A(new_n283_), .ZN(new_n484_));
  NOR3_X1   g347(.A1(new_n459_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g348(.A1(new_n467_), .A2(new_n283_), .ZN(new_n486_));
  AOI21_X1  g349(.A(new_n485_), .B1(new_n486_), .B2(new_n483_), .ZN(G1327gat));
  INV_X1    g350(.A(new_n457_), .ZN(new_n488_));
  NOR2_X1   g351(.A1(new_n488_), .A2(new_n440_), .ZN(new_n489_));
  INV_X1    g352(.A(KEYINPUT40), .ZN(new_n490_));
  AOI21_X1  g353(.A(new_n490_), .B1(new_n336_), .B2(new_n379_), .ZN(new_n491_));
  INV_X1    g354(.A(new_n304_), .ZN(new_n492_));
  OAI21_X1  g355(.A(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n493_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n494_));
  NAND2_X1  g357(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g358(.A(new_n492_), .B1(new_n495_), .B2(new_n334_), .ZN(new_n496_));
  NOR3_X1   g359(.A1(new_n496_), .A2(KEYINPUT40), .A3(new_n380_), .ZN(new_n497_));
  OAI211_X1 g360(.A(new_n251_), .B(new_n489_), .C1(new_n491_), .C2(new_n497_), .ZN(new_n498_));
  AND3_X1   g361(.A1(new_n498_), .A2(KEYINPUT41), .A3(G29gat), .ZN(new_n499_));
  AOI21_X1  g362(.A(KEYINPUT41), .B1(new_n498_), .B2(G29gat), .ZN(new_n500_));
  INV_X1    g363(.A(new_n439_), .ZN(new_n501_));
  NOR2_X1   g364(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g365(.A1(new_n488_), .A2(new_n380_), .ZN(new_n503_));
  NAND2_X1  g366(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g367(.A(KEYINPUT42), .ZN(new_n505_));
  NAND2_X1  g368(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g369(.A1(new_n502_), .A2(KEYINPUT42), .A3(new_n503_), .ZN(new_n507_));
  NAND3_X1  g370(.A1(new_n506_), .A2(new_n416_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g371(.A1(new_n251_), .A2(new_n360_), .ZN(new_n509_));
  OAI22_X1  g372(.A1(new_n499_), .A2(new_n500_), .B1(new_n508_), .B2(new_n509_), .ZN(G1328gat));
  INV_X1    g373(.A(new_n489_), .ZN(new_n511_));
  NAND3_X1  g374(.A1(new_n336_), .A2(new_n490_), .A3(new_n379_), .ZN(new_n512_));
  OAI21_X1  g375(.A(KEYINPUT40), .B1(new_n496_), .B2(new_n380_), .ZN(new_n513_));
  AOI21_X1  g376(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AND2_X1   g377(.A1(new_n514_), .A2(new_n302_), .ZN(new_n515_));
  INV_X1    g378(.A(G36gat), .ZN(new_n516_));
  OAI21_X1  g379(.A(new_n516_), .B1(new_n323_), .B2(KEYINPUT43), .ZN(new_n517_));
  OAI21_X1  g380(.A(new_n517_), .B1(KEYINPUT43), .B2(new_n516_), .ZN(new_n518_));
  OAI22_X1  g381(.A1(new_n515_), .A2(new_n516_), .B1(new_n508_), .B2(new_n518_), .ZN(G1329gat));
  NAND4_X1  g382(.A1(new_n506_), .A2(new_n206_), .A3(new_n416_), .A4(new_n507_), .ZN(new_n520_));
  INV_X1    g383(.A(G43gat), .ZN(new_n521_));
  NOR2_X1   g384(.A1(new_n330_), .A2(new_n521_), .ZN(new_n522_));
  AOI22_X1  g385(.A1(new_n520_), .A2(new_n521_), .B1(new_n514_), .B2(new_n522_), .ZN(G1330gat));
  NAND4_X1  g386(.A1(new_n506_), .A2(new_n283_), .A3(new_n416_), .A4(new_n507_), .ZN(new_n524_));
  INV_X1    g387(.A(G50gat), .ZN(new_n525_));
  NOR2_X1   g388(.A1(new_n484_), .A2(new_n525_), .ZN(new_n526_));
  AOI22_X1  g389(.A1(new_n524_), .A2(new_n525_), .B1(new_n514_), .B2(new_n526_), .ZN(G1331gat));
  NOR2_X1   g390(.A1(new_n416_), .A2(new_n439_), .ZN(new_n528_));
  INV_X1    g391(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g392(.A1(new_n529_), .A2(new_n457_), .ZN(new_n530_));
  NAND3_X1  g393(.A1(new_n336_), .A2(new_n380_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g394(.A(G57gat), .ZN(new_n532_));
  NOR3_X1   g395(.A1(new_n531_), .A2(new_n532_), .A3(new_n252_), .ZN(new_n533_));
  NOR2_X1   g396(.A1(new_n496_), .A2(new_n529_), .ZN(new_n534_));
  NAND3_X1  g397(.A1(new_n534_), .A2(new_n251_), .A3(new_n462_), .ZN(new_n535_));
  AOI21_X1  g398(.A(new_n533_), .B1(new_n532_), .B2(new_n535_), .ZN(G1332gat));
  NAND2_X1  g399(.A1(new_n534_), .A2(new_n462_), .ZN(new_n537_));
  OR3_X1    g400(.A1(new_n537_), .A2(G64gat), .A3(new_n323_), .ZN(new_n538_));
  OR2_X1    g401(.A1(new_n531_), .A2(new_n323_), .ZN(new_n539_));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n540_));
  AND3_X1   g403(.A1(new_n539_), .A2(new_n540_), .A3(G64gat), .ZN(new_n541_));
  AOI21_X1  g404(.A(new_n540_), .B1(new_n539_), .B2(G64gat), .ZN(new_n542_));
  OAI21_X1  g405(.A(new_n538_), .B1(new_n541_), .B2(new_n542_), .ZN(G1333gat));
  NOR2_X1   g406(.A1(new_n531_), .A2(new_n330_), .ZN(new_n544_));
  XNOR2_X1  g407(.A(KEYINPUT10), .B(G71gat), .ZN(new_n545_));
  OR2_X1    g408(.A1(new_n474_), .A2(new_n545_), .ZN(new_n546_));
  OAI22_X1  g409(.A1(new_n544_), .A2(new_n384_), .B1(new_n537_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g410(.A(KEYINPUT45), .ZN(new_n548_));
  XNOR2_X1  g411(.A(new_n547_), .B(new_n548_), .ZN(G1334gat));
  OAI21_X1  g412(.A(G78gat), .B1(new_n531_), .B2(new_n484_), .ZN(new_n550_));
  NAND2_X1  g413(.A1(new_n283_), .A2(new_n382_), .ZN(new_n551_));
  OAI21_X1  g414(.A(new_n550_), .B1(new_n537_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g415(.A(KEYINPUT46), .ZN(new_n553_));
  XNOR2_X1  g416(.A(new_n552_), .B(new_n553_), .ZN(G1335gat));
  NOR2_X1   g417(.A1(new_n529_), .A2(new_n488_), .ZN(new_n555_));
  INV_X1    g418(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g419(.A(new_n556_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n557_));
  NOR2_X1   g420(.A1(new_n252_), .A2(new_n342_), .ZN(new_n558_));
  NAND3_X1  g421(.A1(new_n534_), .A2(new_n251_), .A3(new_n503_), .ZN(new_n559_));
  AOI22_X1  g422(.A1(new_n557_), .A2(new_n558_), .B1(new_n342_), .B2(new_n559_), .ZN(G1336gat));
  OAI211_X1 g423(.A(new_n302_), .B(new_n555_), .C1(new_n491_), .C2(new_n497_), .ZN(new_n561_));
  AND3_X1   g424(.A1(new_n561_), .A2(KEYINPUT47), .A3(G92gat), .ZN(new_n562_));
  AOI21_X1  g425(.A(KEYINPUT47), .B1(new_n561_), .B2(G92gat), .ZN(new_n563_));
  NAND2_X1  g426(.A1(new_n534_), .A2(new_n503_), .ZN(new_n564_));
  NAND2_X1  g427(.A1(new_n302_), .A2(new_n343_), .ZN(new_n565_));
  OAI22_X1  g428(.A1(new_n562_), .A2(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(G1337gat));
  INV_X1    g429(.A(new_n557_), .ZN(new_n567_));
  OAI211_X1 g430(.A(KEYINPUT48), .B(G99gat), .C1(new_n567_), .C2(new_n330_), .ZN(new_n568_));
  INV_X1    g431(.A(KEYINPUT48), .ZN(new_n569_));
  AOI211_X1 g432(.A(new_n330_), .B(new_n556_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n570_));
  INV_X1    g433(.A(G99gat), .ZN(new_n571_));
  OAI21_X1  g434(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g435(.A1(new_n534_), .A2(new_n571_), .A3(new_n206_), .A4(new_n503_), .ZN(new_n573_));
  XNOR2_X1  g436(.A(new_n573_), .B(KEYINPUT49), .ZN(new_n574_));
  NAND3_X1  g437(.A1(new_n568_), .A2(new_n572_), .A3(new_n574_), .ZN(G1338gat));
  INV_X1    g438(.A(G106gat), .ZN(new_n576_));
  AOI21_X1  g439(.A(new_n576_), .B1(new_n557_), .B2(new_n283_), .ZN(new_n577_));
  NAND2_X1  g440(.A1(new_n283_), .A2(new_n576_), .ZN(new_n578_));
  NOR2_X1   g441(.A1(new_n564_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g442(.A(KEYINPUT50), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g443(.A(new_n579_), .ZN(new_n581_));
  INV_X1    g444(.A(KEYINPUT50), .ZN(new_n582_));
  AOI211_X1 g445(.A(new_n484_), .B(new_n556_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n583_));
  OAI211_X1 g446(.A(new_n581_), .B(new_n582_), .C1(new_n583_), .C2(new_n576_), .ZN(new_n584_));
  NAND2_X1  g447(.A1(new_n580_), .A2(new_n584_), .ZN(G1339gat));
  NOR2_X1   g448(.A1(new_n427_), .A2(new_n429_), .ZN(new_n586_));
  NOR2_X1   g449(.A1(new_n426_), .A2(new_n428_), .ZN(new_n587_));
  OAI21_X1  g450(.A(new_n436_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g451(.A1(new_n588_), .A2(new_n438_), .ZN(new_n589_));
  AOI21_X1  g452(.A(new_n589_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n590_));
  NOR2_X1   g453(.A1(new_n590_), .A2(new_n379_), .ZN(new_n591_));
  INV_X1    g454(.A(KEYINPUT52), .ZN(new_n592_));
  NAND2_X1  g455(.A1(new_n401_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g456(.A(new_n395_), .ZN(new_n594_));
  NAND2_X1  g457(.A1(new_n400_), .A2(new_n397_), .ZN(new_n595_));
  OAI21_X1  g458(.A(new_n402_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g459(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g460(.A(new_n592_), .B(new_n402_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n598_));
  NAND2_X1  g461(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g462(.A1(new_n599_), .A2(new_n410_), .ZN(new_n600_));
  INV_X1    g463(.A(KEYINPUT51), .ZN(new_n601_));
  NAND2_X1  g464(.A1(new_n414_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g465(.A1(new_n401_), .A2(KEYINPUT51), .A3(new_n413_), .A4(new_n405_), .ZN(new_n603_));
  AND2_X1   g466(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g467(.A1(new_n600_), .A2(new_n604_), .A3(new_n439_), .ZN(new_n605_));
  AOI21_X1  g468(.A(new_n488_), .B1(new_n591_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g469(.A(new_n589_), .ZN(new_n607_));
  NAND4_X1  g470(.A1(new_n600_), .A2(new_n604_), .A3(KEYINPUT53), .A4(new_n607_), .ZN(new_n608_));
  INV_X1    g471(.A(KEYINPUT53), .ZN(new_n609_));
  NAND4_X1  g472(.A1(new_n602_), .A2(new_n438_), .A3(new_n588_), .A4(new_n603_), .ZN(new_n610_));
  INV_X1    g473(.A(new_n410_), .ZN(new_n611_));
  AOI21_X1  g474(.A(new_n611_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n612_));
  OAI21_X1  g475(.A(new_n609_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g476(.A1(new_n608_), .A2(new_n379_), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g477(.A1(new_n439_), .A2(new_n415_), .ZN(new_n615_));
  AOI22_X1  g478(.A1(new_n606_), .A2(new_n614_), .B1(new_n462_), .B2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g479(.A1(new_n616_), .A2(new_n474_), .A3(new_n283_), .ZN(new_n617_));
  NOR2_X1   g480(.A1(new_n252_), .A2(new_n302_), .ZN(new_n618_));
  NAND2_X1  g481(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g482(.A1(new_n619_), .A2(new_n501_), .ZN(new_n620_));
  XOR2_X1   g483(.A(KEYINPUT54), .B(G113gat), .Z(new_n621_));
  XNOR2_X1  g484(.A(new_n620_), .B(new_n621_), .ZN(G1340gat));
  OAI22_X1  g485(.A1(new_n619_), .A2(new_n416_), .B1(KEYINPUT55), .B2(G120gat), .ZN(new_n623_));
  NAND2_X1  g486(.A1(KEYINPUT55), .A2(G120gat), .ZN(new_n624_));
  XNOR2_X1  g487(.A(new_n623_), .B(new_n624_), .ZN(G1341gat));
  NOR2_X1   g488(.A1(new_n619_), .A2(new_n457_), .ZN(new_n626_));
  XNOR2_X1  g489(.A(new_n626_), .B(new_n168_), .ZN(G1342gat));
  NOR3_X1   g490(.A1(new_n380_), .A2(new_n252_), .A3(new_n302_), .ZN(new_n628_));
  NAND2_X1  g491(.A1(new_n617_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g492(.A(new_n629_), .B(G134gat), .ZN(G1343gat));
  NAND2_X1  g493(.A1(new_n330_), .A2(new_n283_), .ZN(new_n631_));
  NAND2_X1  g494(.A1(new_n606_), .A2(new_n614_), .ZN(new_n632_));
  NAND2_X1  g495(.A1(new_n462_), .A2(new_n615_), .ZN(new_n633_));
  AOI21_X1  g496(.A(new_n631_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AND2_X1   g497(.A1(new_n634_), .A2(new_n618_), .ZN(new_n635_));
  NAND2_X1  g498(.A1(new_n635_), .A2(new_n439_), .ZN(new_n636_));
  XNOR2_X1  g499(.A(new_n636_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g500(.A1(new_n635_), .A2(new_n415_), .ZN(new_n638_));
  XNOR2_X1  g501(.A(new_n638_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g502(.A1(new_n635_), .A2(new_n488_), .ZN(new_n640_));
  XNOR2_X1  g503(.A(new_n640_), .B(G155gat), .ZN(G1346gat));
  NAND2_X1  g504(.A1(new_n634_), .A2(new_n628_), .ZN(new_n642_));
  XNOR2_X1  g505(.A(new_n642_), .B(G162gat), .ZN(G1347gat));
  INV_X1    g506(.A(new_n614_), .ZN(new_n644_));
  AND3_X1   g507(.A1(new_n600_), .A2(new_n604_), .A3(new_n439_), .ZN(new_n645_));
  OAI211_X1 g508(.A(new_n378_), .B(new_n374_), .C1(new_n416_), .C2(new_n589_), .ZN(new_n646_));
  OAI21_X1  g509(.A(new_n457_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g510(.A(new_n633_), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g511(.A1(new_n206_), .A2(new_n252_), .A3(new_n302_), .ZN(new_n649_));
  INV_X1    g512(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g513(.A1(new_n648_), .A2(new_n484_), .A3(new_n650_), .ZN(new_n651_));
  NOR2_X1   g514(.A1(new_n651_), .A2(new_n501_), .ZN(new_n652_));
  XNOR2_X1  g515(.A(new_n652_), .B(new_n147_), .ZN(G1348gat));
  NOR4_X1   g516(.A1(new_n616_), .A2(new_n283_), .A3(new_n416_), .A4(new_n649_), .ZN(new_n654_));
  AOI21_X1  g517(.A(KEYINPUT57), .B1(new_n654_), .B2(new_n148_), .ZN(new_n655_));
  NAND4_X1  g518(.A1(new_n648_), .A2(new_n484_), .A3(new_n415_), .A4(new_n650_), .ZN(new_n656_));
  INV_X1    g519(.A(KEYINPUT57), .ZN(new_n657_));
  NOR3_X1   g520(.A1(new_n656_), .A2(new_n657_), .A3(G176gat), .ZN(new_n658_));
  INV_X1    g521(.A(KEYINPUT56), .ZN(new_n659_));
  AND3_X1   g522(.A1(new_n656_), .A2(new_n659_), .A3(G176gat), .ZN(new_n660_));
  AOI21_X1  g523(.A(new_n659_), .B1(new_n656_), .B2(G176gat), .ZN(new_n661_));
  OAI22_X1  g524(.A1(new_n655_), .A2(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g525(.A(KEYINPUT58), .ZN(new_n663_));
  NAND2_X1  g526(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g527(.A1(new_n654_), .A2(KEYINPUT57), .A3(new_n148_), .ZN(new_n665_));
  OAI21_X1  g528(.A(new_n657_), .B1(new_n656_), .B2(G176gat), .ZN(new_n666_));
  NAND2_X1  g529(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g530(.A(new_n667_), .B(KEYINPUT58), .C1(new_n661_), .C2(new_n660_), .ZN(new_n668_));
  NAND2_X1  g531(.A1(new_n664_), .A2(new_n668_), .ZN(G1349gat));
  NOR2_X1   g532(.A1(new_n651_), .A2(new_n457_), .ZN(new_n670_));
  XNOR2_X1  g533(.A(new_n670_), .B(new_n143_), .ZN(G1350gat));
  OR2_X1    g534(.A1(new_n651_), .A2(new_n380_), .ZN(new_n672_));
  NAND2_X1  g535(.A1(new_n672_), .A2(G190gat), .ZN(new_n673_));
  INV_X1    g536(.A(KEYINPUT59), .ZN(new_n674_));
  NAND2_X1  g537(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g538(.A1(new_n672_), .A2(KEYINPUT59), .A3(G190gat), .ZN(new_n676_));
  NAND2_X1  g539(.A1(new_n159_), .A2(new_n161_), .ZN(new_n677_));
  OAI211_X1 g540(.A(new_n675_), .B(new_n676_), .C1(new_n677_), .C2(new_n672_), .ZN(G1351gat));
  INV_X1    g541(.A(new_n631_), .ZN(new_n679_));
  NAND4_X1  g542(.A1(new_n648_), .A2(new_n252_), .A3(new_n302_), .A4(new_n679_), .ZN(new_n680_));
  NAND2_X1  g543(.A1(new_n680_), .A2(KEYINPUT60), .ZN(new_n681_));
  INV_X1    g544(.A(KEYINPUT60), .ZN(new_n682_));
  NAND4_X1  g545(.A1(new_n634_), .A2(new_n682_), .A3(new_n252_), .A4(new_n302_), .ZN(new_n683_));
  NAND3_X1  g546(.A1(new_n681_), .A2(new_n439_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g547(.A1(new_n684_), .A2(G197gat), .ZN(new_n685_));
  NOR3_X1   g548(.A1(new_n616_), .A2(new_n251_), .A3(new_n631_), .ZN(new_n686_));
  OR2_X1    g549(.A1(new_n686_), .A2(KEYINPUT61), .ZN(new_n687_));
  NAND2_X1  g550(.A1(new_n686_), .A2(KEYINPUT61), .ZN(new_n688_));
  NAND3_X1  g551(.A1(new_n687_), .A2(new_n302_), .A3(new_n688_), .ZN(new_n689_));
  OR2_X1    g552(.A1(new_n501_), .A2(G197gat), .ZN(new_n690_));
  OAI21_X1  g553(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(G1352gat));
  NAND3_X1  g554(.A1(new_n681_), .A2(new_n415_), .A3(new_n683_), .ZN(new_n692_));
  AND3_X1   g555(.A1(new_n692_), .A2(KEYINPUT62), .A3(G204gat), .ZN(new_n693_));
  AOI21_X1  g556(.A(KEYINPUT62), .B1(new_n692_), .B2(G204gat), .ZN(new_n694_));
  OR2_X1    g557(.A1(new_n416_), .A2(G204gat), .ZN(new_n695_));
  OAI22_X1  g558(.A1(new_n693_), .A2(new_n694_), .B1(new_n689_), .B2(new_n695_), .ZN(G1353gat));
  NAND3_X1  g559(.A1(new_n681_), .A2(new_n488_), .A3(new_n683_), .ZN(new_n697_));
  AND3_X1   g560(.A1(new_n697_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n698_));
  AOI21_X1  g561(.A(KEYINPUT63), .B1(new_n697_), .B2(G211gat), .ZN(new_n699_));
  NAND2_X1  g562(.A1(new_n488_), .A2(new_n253_), .ZN(new_n700_));
  OAI22_X1  g563(.A1(new_n698_), .A2(new_n699_), .B1(new_n689_), .B2(new_n700_), .ZN(G1354gat));
  NAND3_X1  g564(.A1(new_n379_), .A2(new_n262_), .A3(new_n264_), .ZN(new_n702_));
  AND3_X1   g565(.A1(new_n681_), .A2(new_n379_), .A3(new_n683_), .ZN(new_n703_));
  OAI22_X1  g566(.A1(new_n689_), .A2(new_n702_), .B1(new_n703_), .B2(new_n254_), .ZN(G1355gat));
endmodule


