//Secret key is'1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_c1908" written by ABC on Wed Nov 16 09:20:44 2022

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G101, G104, G107, G110, G113, G116, G119,
    G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217,
    G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902,
    G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G101, G104, G107, G110, G113,
    G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210,
    G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898,
    G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187_));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188_));
  XNOR2_X1  g002(.A(new_n188_), .B(KEYINPUT22), .ZN(new_n189_));
  INV_X1    g003(.A(new_n189_), .ZN(new_n190_));
  OR2_X1    g004(.A1(KEYINPUT7), .A2(G104), .ZN(new_n191_));
  NAND2_X1  g005(.A1(KEYINPUT7), .A2(G104), .ZN(new_n192_));
  NAND3_X1  g006(.A1(new_n191_), .A2(G107), .A3(new_n192_), .ZN(new_n193_));
  INV_X1    g007(.A(G101), .ZN(new_n194_));
  INV_X1    g008(.A(G107), .ZN(new_n195_));
  NAND3_X1  g009(.A1(new_n195_), .A2(KEYINPUT6), .A3(G104), .ZN(new_n196_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n197_));
  INV_X1    g011(.A(G104), .ZN(new_n198_));
  OAI21_X1  g012(.A(new_n197_), .B1(new_n198_), .B2(G107), .ZN(new_n199_));
  NAND4_X1  g013(.A1(new_n193_), .A2(new_n194_), .A3(new_n196_), .A4(new_n199_), .ZN(new_n200_));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n201_));
  NAND2_X1  g015(.A1(new_n200_), .A2(new_n201_), .ZN(new_n202_));
  AND2_X1   g016(.A1(new_n199_), .A2(new_n196_), .ZN(new_n203_));
  NAND4_X1  g017(.A1(new_n203_), .A2(KEYINPUT9), .A3(new_n194_), .A4(new_n193_), .ZN(new_n204_));
  AND2_X1   g018(.A1(new_n202_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g019(.A(G113), .ZN(new_n206_));
  INV_X1    g020(.A(G119), .ZN(new_n207_));
  NAND2_X1  g021(.A1(new_n207_), .A2(G116), .ZN(new_n208_));
  INV_X1    g022(.A(G116), .ZN(new_n209_));
  NAND2_X1  g023(.A1(new_n209_), .A2(G119), .ZN(new_n210_));
  AOI21_X1  g024(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g025(.A1(new_n211_), .A2(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g026(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g027(.A1(new_n208_), .A2(KEYINPUT4), .ZN(new_n214_));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n215_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n207_), .A3(G116), .ZN(new_n216_));
  NAND4_X1  g030(.A1(new_n214_), .A2(new_n216_), .A3(new_n206_), .A4(new_n210_), .ZN(new_n217_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n218_));
  AOI211_X1 g032(.A(new_n218_), .B(new_n206_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n219_));
  INV_X1    g033(.A(new_n219_), .ZN(new_n220_));
  AND3_X1   g034(.A1(new_n213_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  AND2_X1   g035(.A1(KEYINPUT7), .A2(G104), .ZN(new_n222_));
  NOR2_X1   g036(.A1(KEYINPUT7), .A2(G104), .ZN(new_n223_));
  OAI21_X1  g037(.A(new_n195_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225_));
  NAND2_X1  g039(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g040(.A(KEYINPUT10), .B(new_n195_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n227_));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228_));
  AOI21_X1  g042(.A(new_n228_), .B1(new_n198_), .B2(G107), .ZN(new_n229_));
  NOR3_X1   g043(.A1(new_n195_), .A2(KEYINPUT11), .A3(G104), .ZN(new_n230_));
  NOR2_X1   g044(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g045(.A1(new_n226_), .A2(new_n227_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n233_));
  AND3_X1   g047(.A1(new_n232_), .A2(new_n233_), .A3(G101), .ZN(new_n234_));
  AOI21_X1  g048(.A(new_n233_), .B1(new_n232_), .B2(G101), .ZN(new_n235_));
  OAI211_X1 g049(.A(new_n205_), .B(new_n221_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g050(.A(KEYINPUT13), .ZN(new_n237_));
  NAND2_X1  g051(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239_));
  XOR2_X1   g053(.A(new_n239_), .B(KEYINPUT3), .Z(new_n240_));
  INV_X1    g054(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g055(.A1(new_n232_), .A2(G101), .ZN(new_n242_));
  NAND2_X1  g056(.A1(new_n242_), .A2(KEYINPUT12), .ZN(new_n243_));
  NAND3_X1  g057(.A1(new_n232_), .A2(new_n233_), .A3(G101), .ZN(new_n244_));
  NAND2_X1  g058(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g059(.A1(new_n212_), .A2(new_n219_), .ZN(new_n246_));
  NAND4_X1  g060(.A1(new_n246_), .A2(new_n202_), .A3(new_n217_), .A4(new_n204_), .ZN(new_n247_));
  INV_X1    g061(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g062(.A1(new_n245_), .A2(KEYINPUT13), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n250_));
  OR2_X1    g064(.A1(new_n217_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g065(.A1(new_n214_), .A2(new_n216_), .A3(new_n210_), .ZN(new_n252_));
  NAND2_X1  g066(.A1(new_n252_), .A2(G113), .ZN(new_n253_));
  NAND2_X1  g067(.A1(new_n217_), .A2(new_n250_), .ZN(new_n254_));
  NAND3_X1  g068(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g069(.A1(new_n203_), .A2(new_n193_), .ZN(new_n256_));
  NAND2_X1  g070(.A1(new_n256_), .A2(G101), .ZN(new_n257_));
  NAND2_X1  g071(.A1(new_n257_), .A2(new_n200_), .ZN(new_n258_));
  AND2_X1   g072(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g073(.A(new_n259_), .ZN(new_n260_));
  NAND4_X1  g074(.A1(new_n238_), .A2(new_n241_), .A3(new_n249_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g075(.A(G143), .ZN(new_n262_));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n262_), .B2(G146), .ZN(new_n263_));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264_));
  INV_X1    g078(.A(G146), .ZN(new_n265_));
  NAND3_X1  g079(.A1(new_n264_), .A2(new_n265_), .A3(G143), .ZN(new_n266_));
  NAND2_X1  g080(.A1(new_n262_), .A2(G146), .ZN(new_n267_));
  NAND3_X1  g081(.A1(new_n263_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g082(.A1(new_n268_), .A2(G128), .ZN(new_n269_));
  INV_X1    g083(.A(G128), .ZN(new_n270_));
  NAND4_X1  g084(.A1(new_n263_), .A2(new_n266_), .A3(new_n270_), .A4(new_n267_), .ZN(new_n271_));
  NAND2_X1  g085(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g086(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g087(.A1(new_n273_), .A2(G125), .ZN(new_n274_));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n275_));
  OR2_X1    g089(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g090(.A1(new_n271_), .A2(new_n275_), .ZN(new_n277_));
  NAND2_X1  g091(.A1(new_n265_), .A2(G143), .ZN(new_n278_));
  NAND2_X1  g092(.A1(new_n267_), .A2(new_n278_), .ZN(new_n279_));
  AOI22_X1  g093(.A1(new_n276_), .A2(new_n277_), .B1(G128), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g094(.A(new_n274_), .B1(new_n280_), .B2(G125), .ZN(new_n281_));
  INV_X1    g095(.A(G953), .ZN(new_n282_));
  AOI21_X1  g096(.A(KEYINPUT16), .B1(new_n282_), .B2(G224), .ZN(new_n283_));
  NAND2_X1  g097(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g098(.A1(new_n281_), .A2(new_n283_), .ZN(new_n285_));
  AOI22_X1  g099(.A1(new_n261_), .A2(KEYINPUT17), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g100(.A(KEYINPUT19), .ZN(new_n287_));
  NAND2_X1  g101(.A1(new_n202_), .A2(new_n204_), .ZN(new_n288_));
  AOI21_X1  g102(.A(new_n288_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n289_));
  OAI21_X1  g103(.A(new_n287_), .B1(new_n289_), .B2(new_n221_), .ZN(new_n290_));
  OAI21_X1  g104(.A(new_n205_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n291_));
  NAND3_X1  g105(.A1(new_n213_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n292_));
  NAND3_X1  g106(.A1(new_n291_), .A2(KEYINPUT19), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g107(.A(new_n247_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n294_));
  NAND2_X1  g108(.A1(new_n294_), .A2(KEYINPUT20), .ZN(new_n295_));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n296_));
  NAND2_X1  g110(.A1(new_n236_), .A2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g111(.A1(new_n290_), .A2(new_n293_), .A3(new_n295_), .A4(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g112(.A(new_n240_), .B(KEYINPUT18), .ZN(new_n299_));
  NAND2_X1  g113(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g114(.A(new_n259_), .B1(new_n294_), .B2(KEYINPUT13), .ZN(new_n301_));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n302_));
  NAND4_X1  g116(.A1(new_n301_), .A2(new_n302_), .A3(new_n241_), .A4(new_n238_), .ZN(new_n303_));
  NAND3_X1  g117(.A1(new_n286_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n305_));
  NAND2_X1  g119(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g120(.A1(new_n286_), .A2(new_n300_), .A3(KEYINPUT21), .A4(new_n303_), .ZN(new_n307_));
  NAND2_X1  g121(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g122(.A(KEYINPUT0), .B(G902), .Z(new_n309_));
  INV_X1    g123(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g124(.A1(new_n261_), .A2(KEYINPUT14), .ZN(new_n311_));
  INV_X1    g125(.A(KEYINPUT14), .ZN(new_n312_));
  NAND4_X1  g126(.A1(new_n301_), .A2(new_n312_), .A3(new_n241_), .A4(new_n238_), .ZN(new_n313_));
  INV_X1    g127(.A(KEYINPUT15), .ZN(new_n314_));
  AOI211_X1 g128(.A(new_n314_), .B(new_n241_), .C1(new_n301_), .C2(new_n238_), .ZN(new_n315_));
  NAND3_X1  g129(.A1(new_n238_), .A2(new_n260_), .A3(new_n249_), .ZN(new_n316_));
  AOI21_X1  g130(.A(KEYINPUT15), .B1(new_n316_), .B2(new_n240_), .ZN(new_n317_));
  OAI211_X1 g131(.A(new_n311_), .B(new_n313_), .C1(new_n315_), .C2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g132(.A1(new_n282_), .A2(G224), .ZN(new_n319_));
  XOR2_X1   g133(.A(new_n281_), .B(new_n319_), .Z(new_n320_));
  AOI21_X1  g134(.A(new_n310_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g135(.A1(new_n308_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g136(.A1(new_n322_), .A2(KEYINPUT23), .ZN(new_n323_));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324_));
  NAND3_X1  g138(.A1(new_n308_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g139(.A(new_n190_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g140(.A(new_n324_), .B1(new_n308_), .B2(new_n321_), .ZN(new_n327_));
  NOR2_X1   g141(.A1(new_n327_), .A2(new_n189_), .ZN(new_n328_));
  OAI21_X1  g142(.A(new_n187_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n330_));
  NAND2_X1  g144(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AND3_X1   g145(.A1(new_n308_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n332_));
  OAI21_X1  g146(.A(new_n189_), .B1(new_n332_), .B2(new_n327_), .ZN(new_n333_));
  NAND2_X1  g147(.A1(new_n323_), .A2(new_n190_), .ZN(new_n334_));
  NAND2_X1  g148(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g149(.A1(new_n335_), .A2(KEYINPUT24), .A3(new_n187_), .ZN(new_n336_));
  AND2_X1   g150(.A1(KEYINPUT25), .A2(G953), .ZN(new_n337_));
  NOR2_X1   g151(.A1(KEYINPUT25), .A2(G953), .ZN(new_n338_));
  NOR2_X1   g152(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g153(.A1(new_n339_), .A2(G952), .ZN(new_n340_));
  INV_X1    g154(.A(G234), .ZN(new_n341_));
  INV_X1    g155(.A(G237), .ZN(new_n342_));
  OAI21_X1  g156(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g157(.A(new_n343_), .B(KEYINPUT50), .ZN(new_n344_));
  INV_X1    g158(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g159(.A(G902), .ZN(new_n346_));
  AOI21_X1  g160(.A(new_n346_), .B1(G234), .B2(G237), .ZN(new_n347_));
  INV_X1    g161(.A(G898), .ZN(new_n348_));
  NAND3_X1  g162(.A1(new_n347_), .A2(new_n348_), .A3(G953), .ZN(new_n349_));
  NAND2_X1  g163(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g164(.A(new_n350_), .B(KEYINPUT51), .Z(new_n351_));
  INV_X1    g165(.A(G475), .ZN(new_n352_));
  NAND2_X1  g166(.A1(new_n309_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g167(.A1(new_n191_), .A2(new_n192_), .ZN(new_n354_));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355_));
  XNOR2_X1  g169(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND3_X1  g170(.A1(new_n342_), .A2(new_n282_), .A3(G214), .ZN(new_n357_));
  AOI21_X1  g171(.A(G131), .B1(new_n357_), .B2(new_n262_), .ZN(new_n358_));
  XNOR2_X1  g172(.A(KEYINPUT40), .B(G237), .ZN(new_n359_));
  NAND4_X1  g173(.A1(new_n339_), .A2(new_n359_), .A3(G143), .A4(G214), .ZN(new_n360_));
  AND2_X1   g174(.A1(new_n360_), .A2(KEYINPUT41), .ZN(new_n361_));
  NOR2_X1   g175(.A1(new_n360_), .A2(KEYINPUT41), .ZN(new_n362_));
  OAI21_X1  g176(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g177(.A(KEYINPUT42), .ZN(new_n364_));
  NAND2_X1  g178(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  AND2_X1   g179(.A1(new_n339_), .A2(new_n359_), .ZN(new_n366_));
  INV_X1    g180(.A(KEYINPUT41), .ZN(new_n367_));
  NAND4_X1  g181(.A1(new_n366_), .A2(new_n367_), .A3(G143), .A4(G214), .ZN(new_n368_));
  NAND2_X1  g182(.A1(new_n360_), .A2(KEYINPUT41), .ZN(new_n369_));
  NAND2_X1  g183(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g184(.A1(new_n370_), .A2(KEYINPUT42), .A3(new_n358_), .ZN(new_n371_));
  NAND2_X1  g185(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  AND2_X1   g186(.A1(new_n366_), .A2(G214), .ZN(new_n373_));
  OAI21_X1  g187(.A(new_n370_), .B1(G143), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g188(.A1(new_n374_), .A2(G131), .ZN(new_n375_));
  NAND2_X1  g189(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g190(.A(G125), .B(G140), .ZN(new_n377_));
  OR2_X1    g191(.A1(new_n377_), .A2(new_n265_), .ZN(new_n378_));
  NAND2_X1  g192(.A1(new_n377_), .A2(new_n265_), .ZN(new_n379_));
  NAND2_X1  g193(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g194(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g195(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g196(.A(new_n382_), .B(KEYINPUT49), .Z(new_n383_));
  AOI21_X1  g197(.A(G143), .B1(new_n357_), .B2(KEYINPUT43), .ZN(new_n384_));
  OAI21_X1  g198(.A(new_n384_), .B1(KEYINPUT43), .B2(new_n357_), .ZN(new_n385_));
  OAI211_X1 g199(.A(KEYINPUT44), .B(new_n385_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n386_));
  NAND2_X1  g200(.A1(new_n386_), .A2(G131), .ZN(new_n387_));
  AOI21_X1  g201(.A(KEYINPUT44), .B1(new_n370_), .B2(new_n385_), .ZN(new_n388_));
  NOR2_X1   g202(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g203(.A(KEYINPUT42), .B1(new_n370_), .B2(new_n358_), .ZN(new_n390_));
  INV_X1    g204(.A(new_n358_), .ZN(new_n391_));
  AOI211_X1 g205(.A(new_n364_), .B(new_n391_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n392_));
  OAI21_X1  g206(.A(new_n380_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g207(.A(KEYINPUT45), .ZN(new_n394_));
  NOR3_X1   g208(.A1(new_n389_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g209(.A1(new_n370_), .A2(new_n385_), .ZN(new_n396_));
  INV_X1    g210(.A(KEYINPUT44), .ZN(new_n397_));
  NAND2_X1  g211(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g212(.A1(new_n398_), .A2(G131), .A3(new_n386_), .ZN(new_n399_));
  AOI21_X1  g213(.A(new_n381_), .B1(new_n365_), .B2(new_n371_), .ZN(new_n400_));
  AOI21_X1  g214(.A(KEYINPUT45), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g215(.A1(new_n395_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g216(.A(new_n356_), .B1(new_n383_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g217(.A(new_n394_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n404_));
  NAND3_X1  g218(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT45), .ZN(new_n405_));
  XOR2_X1   g219(.A(new_n380_), .B(KEYINPUT39), .Z(new_n406_));
  INV_X1    g220(.A(new_n406_), .ZN(new_n407_));
  AOI22_X1  g221(.A1(new_n404_), .A2(new_n405_), .B1(new_n376_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g222(.A(new_n356_), .ZN(new_n409_));
  NAND2_X1  g223(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g224(.A(new_n353_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g225(.A1(new_n376_), .A2(new_n407_), .ZN(new_n412_));
  AOI21_X1  g226(.A(KEYINPUT46), .B1(new_n356_), .B2(KEYINPUT47), .ZN(new_n413_));
  OAI211_X1 g227(.A(new_n412_), .B(new_n413_), .C1(new_n395_), .C2(new_n401_), .ZN(new_n414_));
  NAND2_X1  g228(.A1(new_n356_), .A2(KEYINPUT47), .ZN(new_n415_));
  OAI21_X1  g229(.A(new_n414_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g230(.A(KEYINPUT46), .ZN(new_n417_));
  AOI21_X1  g231(.A(new_n417_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n418_));
  OAI21_X1  g232(.A(new_n346_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g233(.A(new_n352_), .B1(new_n419_), .B2(KEYINPUT48), .ZN(new_n420_));
  INV_X1    g234(.A(KEYINPUT48), .ZN(new_n421_));
  OAI211_X1 g235(.A(new_n421_), .B(new_n346_), .C1(new_n416_), .C2(new_n418_), .ZN(new_n422_));
  AOI21_X1  g236(.A(new_n411_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g237(.A(G478), .ZN(new_n424_));
  XNOR2_X1  g238(.A(G116), .B(G122), .ZN(new_n425_));
  XNOR2_X1  g239(.A(new_n425_), .B(G107), .ZN(new_n426_));
  INV_X1    g240(.A(G134), .ZN(new_n427_));
  NAND2_X1  g241(.A1(new_n262_), .A2(G128), .ZN(new_n428_));
  NAND2_X1  g242(.A1(new_n270_), .A2(G143), .ZN(new_n429_));
  AOI21_X1  g243(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g244(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g245(.A1(new_n428_), .A2(KEYINPUT34), .ZN(new_n432_));
  INV_X1    g246(.A(KEYINPUT34), .ZN(new_n433_));
  NAND3_X1  g247(.A1(new_n433_), .A2(new_n262_), .A3(G128), .ZN(new_n434_));
  NAND3_X1  g248(.A1(new_n432_), .A2(new_n434_), .A3(new_n429_), .ZN(new_n435_));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n436_));
  OR3_X1    g250(.A1(new_n435_), .A2(new_n436_), .A3(G134), .ZN(new_n437_));
  OAI21_X1  g251(.A(new_n436_), .B1(new_n435_), .B2(G134), .ZN(new_n438_));
  NAND3_X1  g252(.A1(new_n431_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n440_));
  NAND2_X1  g254(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g255(.A1(new_n431_), .A2(KEYINPUT36), .A3(new_n437_), .A4(new_n438_), .ZN(new_n442_));
  NAND2_X1  g256(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g257(.A1(new_n282_), .A2(G217), .A3(G234), .ZN(new_n444_));
  XNOR2_X1  g258(.A(new_n444_), .B(KEYINPUT33), .ZN(new_n445_));
  XNOR2_X1  g259(.A(new_n435_), .B(G134), .ZN(new_n446_));
  NAND2_X1  g260(.A1(new_n209_), .A2(G122), .ZN(new_n447_));
  AOI21_X1  g261(.A(new_n195_), .B1(new_n447_), .B2(KEYINPUT37), .ZN(new_n448_));
  XNOR2_X1  g262(.A(new_n448_), .B(new_n425_), .ZN(new_n449_));
  NAND2_X1  g263(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g264(.A1(new_n443_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g265(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g266(.A(new_n445_), .B1(new_n443_), .B2(new_n450_), .ZN(new_n453_));
  OAI211_X1 g267(.A(new_n424_), .B(new_n309_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g268(.A1(new_n454_), .A2(KEYINPUT38), .ZN(new_n455_));
  OAI21_X1  g269(.A(new_n309_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n456_));
  NAND2_X1  g270(.A1(new_n456_), .A2(G478), .ZN(new_n457_));
  XNOR2_X1  g271(.A(new_n455_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g272(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g273(.A1(new_n423_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g274(.A(new_n460_), .ZN(new_n461_));
  NAND4_X1  g275(.A1(new_n331_), .A2(new_n336_), .A3(new_n351_), .A4(new_n461_), .ZN(new_n462_));
  OAI21_X1  g276(.A(G221), .B1(new_n341_), .B2(G902), .ZN(new_n463_));
  INV_X1    g277(.A(G469), .ZN(new_n464_));
  NAND2_X1  g278(.A1(new_n309_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g279(.A1(new_n258_), .A2(new_n272_), .ZN(new_n466_));
  INV_X1    g280(.A(new_n466_), .ZN(new_n467_));
  OAI211_X1 g281(.A(new_n280_), .B(new_n205_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n468_));
  INV_X1    g282(.A(new_n468_), .ZN(new_n469_));
  AOI21_X1  g283(.A(new_n467_), .B1(new_n469_), .B2(KEYINPUT26), .ZN(new_n470_));
  INV_X1    g284(.A(G131), .ZN(new_n471_));
  NAND2_X1  g285(.A1(new_n427_), .A2(G137), .ZN(new_n472_));
  INV_X1    g286(.A(G137), .ZN(new_n473_));
  NAND3_X1  g287(.A1(new_n473_), .A2(KEYINPUT27), .A3(G134), .ZN(new_n474_));
  INV_X1    g288(.A(new_n474_), .ZN(new_n475_));
  AOI21_X1  g289(.A(KEYINPUT27), .B1(new_n473_), .B2(G134), .ZN(new_n476_));
  OAI211_X1 g290(.A(new_n471_), .B(new_n472_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g291(.A1(new_n477_), .A2(KEYINPUT28), .ZN(new_n478_));
  NAND2_X1  g292(.A1(new_n473_), .A2(G134), .ZN(new_n479_));
  INV_X1    g293(.A(KEYINPUT27), .ZN(new_n480_));
  NAND2_X1  g294(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g295(.A1(new_n481_), .A2(new_n474_), .ZN(new_n482_));
  INV_X1    g296(.A(KEYINPUT28), .ZN(new_n483_));
  NAND4_X1  g297(.A1(new_n482_), .A2(new_n483_), .A3(new_n471_), .A4(new_n472_), .ZN(new_n484_));
  OAI21_X1  g298(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n485_));
  NAND2_X1  g299(.A1(new_n485_), .A2(G131), .ZN(new_n486_));
  AND3_X1   g300(.A1(new_n478_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g301(.A(KEYINPUT26), .ZN(new_n488_));
  NAND2_X1  g302(.A1(new_n468_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g303(.A1(new_n470_), .A2(KEYINPUT29), .A3(new_n487_), .A4(new_n489_), .ZN(new_n490_));
  NAND4_X1  g304(.A1(new_n245_), .A2(KEYINPUT26), .A3(new_n280_), .A4(new_n205_), .ZN(new_n491_));
  NAND4_X1  g305(.A1(new_n489_), .A2(new_n491_), .A3(new_n487_), .A4(new_n466_), .ZN(new_n492_));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n493_));
  NAND2_X1  g307(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g308(.A1(new_n489_), .A2(new_n491_), .A3(new_n466_), .ZN(new_n495_));
  NAND3_X1  g309(.A1(new_n478_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n496_));
  NAND2_X1  g310(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g311(.A1(new_n490_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g312(.A1(new_n339_), .A2(G227), .ZN(new_n499_));
  XNOR2_X1  g313(.A(G110), .B(G140), .ZN(new_n500_));
  XNOR2_X1  g314(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g315(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g316(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504_));
  OR2_X1    g318(.A1(new_n492_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g319(.A1(new_n289_), .A2(new_n280_), .ZN(new_n506_));
  OAI21_X1  g320(.A(new_n496_), .B1(new_n506_), .B2(new_n469_), .ZN(new_n507_));
  NAND2_X1  g321(.A1(new_n492_), .A2(new_n504_), .ZN(new_n508_));
  NAND4_X1  g322(.A1(new_n505_), .A2(new_n501_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g323(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g324(.A1(new_n510_), .A2(KEYINPUT31), .ZN(new_n511_));
  INV_X1    g325(.A(KEYINPUT31), .ZN(new_n512_));
  NAND3_X1  g326(.A1(new_n503_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g327(.A(new_n465_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g328(.A1(new_n505_), .A2(new_n502_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n515_));
  AND2_X1   g329(.A1(new_n515_), .A2(new_n309_), .ZN(new_n516_));
  NAND2_X1  g330(.A1(new_n498_), .A2(new_n501_), .ZN(new_n517_));
  AOI21_X1  g331(.A(new_n464_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g332(.A(new_n463_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n520_));
  NAND2_X1  g334(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g335(.A(KEYINPUT32), .B(new_n463_), .C1(new_n514_), .C2(new_n518_), .ZN(new_n522_));
  NAND2_X1  g336(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g337(.A1(new_n462_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g338(.A(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n526_));
  NAND2_X1  g340(.A1(new_n279_), .A2(G128), .ZN(new_n527_));
  AND2_X1   g341(.A1(new_n271_), .A2(new_n275_), .ZN(new_n528_));
  NOR2_X1   g342(.A1(new_n271_), .A2(new_n275_), .ZN(new_n529_));
  OAI21_X1  g343(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g344(.A(KEYINPUT58), .B1(new_n473_), .B2(G134), .ZN(new_n531_));
  INV_X1    g345(.A(KEYINPUT58), .ZN(new_n532_));
  NAND3_X1  g346(.A1(new_n532_), .A2(new_n427_), .A3(G137), .ZN(new_n533_));
  NAND3_X1  g347(.A1(new_n531_), .A2(new_n533_), .A3(new_n479_), .ZN(new_n534_));
  NAND2_X1  g348(.A1(new_n534_), .A2(G131), .ZN(new_n535_));
  INV_X1    g349(.A(KEYINPUT59), .ZN(new_n536_));
  NAND2_X1  g350(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g351(.A1(new_n534_), .A2(KEYINPUT59), .A3(G131), .ZN(new_n538_));
  NAND3_X1  g352(.A1(new_n537_), .A2(new_n538_), .A3(new_n477_), .ZN(new_n539_));
  NOR2_X1   g353(.A1(new_n530_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g354(.A(KEYINPUT60), .ZN(new_n541_));
  OAI21_X1  g355(.A(new_n541_), .B1(new_n487_), .B2(new_n273_), .ZN(new_n542_));
  NAND3_X1  g356(.A1(new_n496_), .A2(KEYINPUT60), .A3(new_n272_), .ZN(new_n543_));
  AOI21_X1  g357(.A(new_n540_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g358(.A(new_n255_), .B(KEYINPUT57), .ZN(new_n545_));
  OAI21_X1  g359(.A(KEYINPUT61), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g360(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  OR2_X1    g361(.A1(new_n530_), .A2(new_n539_), .ZN(new_n548_));
  AND3_X1   g362(.A1(new_n496_), .A2(KEYINPUT60), .A3(new_n272_), .ZN(new_n549_));
  AOI21_X1  g363(.A(KEYINPUT60), .B1(new_n496_), .B2(new_n272_), .ZN(new_n550_));
  OAI21_X1  g364(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g365(.A(KEYINPUT61), .ZN(new_n552_));
  INV_X1    g366(.A(KEYINPUT57), .ZN(new_n553_));
  XNOR2_X1  g367(.A(new_n255_), .B(new_n553_), .ZN(new_n554_));
  NAND3_X1  g368(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g369(.A1(new_n546_), .A2(new_n547_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g370(.A(KEYINPUT65), .ZN(new_n557_));
  AND2_X1   g371(.A1(new_n366_), .A2(G210), .ZN(new_n558_));
  XNOR2_X1  g372(.A(KEYINPUT56), .B(G101), .ZN(new_n559_));
  XNOR2_X1  g373(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g374(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g375(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  AND2_X1   g376(.A1(new_n556_), .A2(new_n561_), .ZN(new_n563_));
  INV_X1    g377(.A(KEYINPUT63), .ZN(new_n564_));
  OAI21_X1  g378(.A(new_n545_), .B1(new_n544_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g379(.A1(new_n551_), .A2(KEYINPUT63), .A3(new_n554_), .ZN(new_n566_));
  NAND3_X1  g380(.A1(new_n565_), .A2(new_n560_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g381(.A1(new_n567_), .A2(KEYINPUT65), .ZN(new_n568_));
  OAI211_X1 g382(.A(new_n309_), .B(new_n562_), .C1(new_n563_), .C2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g383(.A(new_n526_), .B1(new_n569_), .B2(G472), .ZN(new_n570_));
  AND3_X1   g384(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n571_));
  NAND2_X1  g385(.A1(new_n556_), .A2(new_n561_), .ZN(new_n572_));
  INV_X1    g386(.A(new_n568_), .ZN(new_n573_));
  AOI21_X1  g387(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g388(.A(G472), .ZN(new_n575_));
  NAND4_X1  g389(.A1(new_n574_), .A2(KEYINPUT66), .A3(new_n575_), .A4(new_n309_), .ZN(new_n576_));
  AND3_X1   g390(.A1(new_n551_), .A2(KEYINPUT63), .A3(new_n554_), .ZN(new_n577_));
  AOI21_X1  g391(.A(new_n554_), .B1(new_n551_), .B2(KEYINPUT63), .ZN(new_n578_));
  OAI21_X1  g392(.A(new_n561_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g393(.A1(new_n546_), .A2(new_n547_), .A3(new_n555_), .A4(new_n560_), .ZN(new_n580_));
  AND3_X1   g394(.A1(new_n579_), .A2(new_n580_), .A3(KEYINPUT62), .ZN(new_n581_));
  NOR2_X1   g395(.A1(new_n580_), .A2(KEYINPUT62), .ZN(new_n582_));
  OAI21_X1  g396(.A(G472), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g397(.A1(new_n309_), .A2(new_n575_), .ZN(new_n584_));
  INV_X1    g398(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g399(.A1(new_n583_), .A2(KEYINPUT64), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g400(.A(KEYINPUT64), .ZN(new_n587_));
  NAND3_X1  g401(.A1(new_n579_), .A2(new_n580_), .A3(KEYINPUT62), .ZN(new_n588_));
  OAI21_X1  g402(.A(new_n588_), .B1(KEYINPUT62), .B2(new_n580_), .ZN(new_n589_));
  OAI211_X1 g403(.A(new_n587_), .B(G472), .C1(new_n589_), .C2(new_n310_), .ZN(new_n590_));
  AOI22_X1  g404(.A1(new_n570_), .A2(new_n576_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g405(.A(KEYINPUT53), .B(G110), .Z(new_n592_));
  XNOR2_X1  g406(.A(G119), .B(G128), .ZN(new_n593_));
  NAND2_X1  g407(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g408(.A(G110), .ZN(new_n595_));
  OAI211_X1 g409(.A(new_n380_), .B(new_n594_), .C1(new_n595_), .C2(new_n593_), .ZN(new_n596_));
  INV_X1    g410(.A(KEYINPUT52), .ZN(new_n597_));
  XNOR2_X1  g411(.A(new_n378_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g412(.A1(new_n593_), .A2(G110), .ZN(new_n599_));
  INV_X1    g413(.A(new_n592_), .ZN(new_n600_));
  OAI211_X1 g414(.A(new_n379_), .B(new_n599_), .C1(new_n600_), .C2(new_n593_), .ZN(new_n601_));
  OAI21_X1  g415(.A(new_n596_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g416(.A1(new_n339_), .A2(G221), .A3(G234), .ZN(new_n603_));
  XNOR2_X1  g417(.A(new_n603_), .B(new_n473_), .ZN(new_n604_));
  NAND2_X1  g418(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g419(.A1(new_n605_), .A2(KEYINPUT54), .ZN(new_n606_));
  OR2_X1    g420(.A1(new_n602_), .A2(new_n604_), .ZN(new_n607_));
  XNOR2_X1  g421(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  AOI21_X1  g422(.A(KEYINPUT55), .B1(new_n608_), .B2(new_n309_), .ZN(new_n609_));
  OAI21_X1  g423(.A(G217), .B1(new_n310_), .B2(new_n341_), .ZN(new_n610_));
  NOR2_X1   g424(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g425(.A1(new_n608_), .A2(KEYINPUT55), .A3(new_n309_), .ZN(new_n612_));
  NAND2_X1  g426(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g427(.A1(new_n608_), .A2(new_n309_), .A3(new_n610_), .ZN(new_n614_));
  NAND2_X1  g428(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g429(.A(new_n525_), .B1(new_n591_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g430(.A1(new_n576_), .A2(new_n570_), .ZN(new_n617_));
  NAND2_X1  g431(.A1(new_n586_), .A2(new_n590_), .ZN(new_n618_));
  NAND2_X1  g432(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g433(.A(new_n615_), .ZN(new_n620_));
  NAND3_X1  g434(.A1(new_n619_), .A2(KEYINPUT67), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g435(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g436(.A1(new_n524_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g437(.A(new_n623_), .B(G101), .ZN(G3));
  NAND3_X1  g438(.A1(new_n572_), .A2(KEYINPUT65), .A3(new_n567_), .ZN(new_n625_));
  NOR2_X1   g439(.A1(G472), .A2(G902), .ZN(new_n626_));
  NAND3_X1  g440(.A1(new_n625_), .A2(new_n562_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g441(.A(KEYINPUT73), .ZN(new_n628_));
  NAND2_X1  g442(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g443(.A1(new_n625_), .A2(KEYINPUT73), .A3(new_n562_), .A4(new_n626_), .ZN(new_n630_));
  NAND2_X1  g444(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g445(.A1(new_n569_), .A2(G472), .ZN(new_n632_));
  NAND2_X1  g446(.A1(new_n632_), .A2(KEYINPUT72), .ZN(new_n633_));
  INV_X1    g447(.A(KEYINPUT72), .ZN(new_n634_));
  NAND3_X1  g448(.A1(new_n569_), .A2(new_n634_), .A3(G472), .ZN(new_n635_));
  NAND3_X1  g449(.A1(new_n631_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  NOR3_X1   g450(.A1(new_n523_), .A2(new_n615_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g451(.A(KEYINPUT24), .B1(new_n335_), .B2(new_n187_), .ZN(new_n638_));
  INV_X1    g452(.A(new_n187_), .ZN(new_n639_));
  AOI211_X1 g453(.A(new_n330_), .B(new_n639_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n640_));
  NOR2_X1   g454(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g455(.A1(new_n443_), .A2(new_n450_), .ZN(new_n642_));
  INV_X1    g456(.A(KEYINPUT69), .ZN(new_n643_));
  XNOR2_X1  g457(.A(new_n445_), .B(KEYINPUT68), .ZN(new_n644_));
  INV_X1    g458(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g459(.A1(new_n642_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g460(.A1(new_n451_), .A2(KEYINPUT69), .ZN(new_n647_));
  AOI21_X1  g461(.A(new_n644_), .B1(new_n443_), .B2(new_n450_), .ZN(new_n648_));
  OAI211_X1 g462(.A(new_n309_), .B(new_n646_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g463(.A1(new_n649_), .A2(G478), .ZN(new_n650_));
  NAND2_X1  g464(.A1(new_n650_), .A2(KEYINPUT70), .ZN(new_n651_));
  INV_X1    g465(.A(KEYINPUT70), .ZN(new_n652_));
  NAND3_X1  g466(.A1(new_n649_), .A2(new_n652_), .A3(G478), .ZN(new_n653_));
  AND4_X1   g467(.A1(KEYINPUT71), .A2(new_n651_), .A3(new_n454_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g468(.A(new_n454_), .ZN(new_n655_));
  AOI21_X1  g469(.A(new_n655_), .B1(new_n650_), .B2(KEYINPUT70), .ZN(new_n656_));
  AOI21_X1  g470(.A(KEYINPUT71), .B1(new_n656_), .B2(new_n653_), .ZN(new_n657_));
  NOR2_X1   g471(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g472(.A1(new_n423_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g473(.A1(new_n637_), .A2(new_n641_), .A3(new_n350_), .A4(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g474(.A(new_n660_), .B(G104), .ZN(G6));
  INV_X1    g475(.A(new_n410_), .ZN(new_n662_));
  NOR2_X1   g476(.A1(new_n408_), .A2(new_n409_), .ZN(new_n663_));
  OAI21_X1  g477(.A(new_n309_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g478(.A(new_n411_), .B1(new_n664_), .B2(G475), .ZN(new_n665_));
  NAND2_X1  g479(.A1(new_n665_), .A2(new_n458_), .ZN(new_n666_));
  INV_X1    g480(.A(new_n666_), .ZN(new_n667_));
  NAND4_X1  g481(.A1(new_n637_), .A2(new_n641_), .A3(new_n350_), .A4(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g482(.A(new_n668_), .B(G107), .ZN(G9));
  INV_X1    g483(.A(KEYINPUT74), .ZN(new_n670_));
  NAND2_X1  g484(.A1(new_n607_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g485(.A(new_n671_), .B(new_n605_), .ZN(new_n672_));
  NAND2_X1  g486(.A1(new_n672_), .A2(new_n610_), .ZN(new_n673_));
  NAND2_X1  g487(.A1(new_n673_), .A2(KEYINPUT75), .ZN(new_n674_));
  INV_X1    g488(.A(KEYINPUT75), .ZN(new_n675_));
  NAND3_X1  g489(.A1(new_n672_), .A2(new_n675_), .A3(new_n610_), .ZN(new_n676_));
  NAND3_X1  g490(.A1(new_n674_), .A2(new_n309_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g491(.A1(new_n677_), .A2(new_n613_), .ZN(new_n678_));
  NAND4_X1  g492(.A1(new_n631_), .A2(new_n633_), .A3(new_n635_), .A4(new_n678_), .ZN(new_n679_));
  INV_X1    g493(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g494(.A1(new_n524_), .A2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g495(.A(KEYINPUT76), .B(G110), .Z(new_n682_));
  XNOR2_X1  g496(.A(new_n681_), .B(new_n682_), .ZN(G12));
  XOR2_X1   g497(.A(KEYINPUT77), .B(G900), .Z(new_n684_));
  NAND3_X1  g498(.A1(new_n684_), .A2(G953), .A3(new_n347_), .ZN(new_n685_));
  XOR2_X1   g499(.A(new_n685_), .B(KEYINPUT78), .Z(new_n686_));
  NOR2_X1   g500(.A1(new_n344_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g501(.A1(new_n666_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g502(.A1(new_n331_), .A2(new_n336_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g503(.A(new_n678_), .ZN(new_n690_));
  AOI21_X1  g504(.A(new_n690_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n691_));
  NAND3_X1  g505(.A1(new_n521_), .A2(new_n522_), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g506(.A(KEYINPUT79), .B1(new_n689_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g507(.A(KEYINPUT79), .ZN(new_n694_));
  AND3_X1   g508(.A1(new_n521_), .A2(new_n522_), .A3(new_n691_), .ZN(new_n695_));
  NAND4_X1  g509(.A1(new_n641_), .A2(new_n694_), .A3(new_n695_), .A4(new_n688_), .ZN(new_n696_));
  NAND2_X1  g510(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g511(.A(KEYINPUT80), .B(G128), .ZN(new_n698_));
  XNOR2_X1  g512(.A(new_n697_), .B(new_n698_), .ZN(G30));
  INV_X1    g513(.A(new_n329_), .ZN(new_n700_));
  OR2_X1    g514(.A1(new_n519_), .A2(new_n687_), .ZN(new_n701_));
  OR2_X1    g515(.A1(new_n701_), .A2(KEYINPUT82), .ZN(new_n702_));
  NAND2_X1  g516(.A1(new_n701_), .A2(KEYINPUT82), .ZN(new_n703_));
  NOR2_X1   g517(.A1(new_n423_), .A2(new_n459_), .ZN(new_n704_));
  INV_X1    g518(.A(new_n567_), .ZN(new_n705_));
  XOR2_X1   g519(.A(new_n547_), .B(KEYINPUT81), .Z(new_n706_));
  NAND3_X1  g520(.A1(new_n706_), .A2(new_n555_), .A3(new_n546_), .ZN(new_n707_));
  AOI21_X1  g521(.A(new_n705_), .B1(new_n707_), .B2(new_n561_), .ZN(new_n708_));
  OAI21_X1  g522(.A(G472), .B1(new_n708_), .B2(G902), .ZN(new_n709_));
  NAND2_X1  g523(.A1(new_n617_), .A2(new_n709_), .ZN(new_n710_));
  AND3_X1   g524(.A1(new_n704_), .A2(new_n690_), .A3(new_n710_), .ZN(new_n711_));
  AND4_X1   g525(.A1(new_n700_), .A2(new_n702_), .A3(new_n703_), .A4(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g526(.A(new_n712_), .B(new_n262_), .ZN(G45));
  NOR3_X1   g527(.A1(new_n423_), .A2(new_n658_), .A3(new_n687_), .ZN(new_n714_));
  NAND4_X1  g528(.A1(new_n695_), .A2(new_n331_), .A3(new_n336_), .A4(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g529(.A(new_n715_), .B(G146), .ZN(G48));
  NAND3_X1  g530(.A1(new_n641_), .A2(new_n350_), .A3(new_n659_), .ZN(new_n717_));
  AND3_X1   g531(.A1(new_n503_), .A2(new_n512_), .A3(new_n509_), .ZN(new_n718_));
  AOI21_X1  g532(.A(new_n512_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n719_));
  OAI211_X1 g533(.A(G469), .B(new_n309_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g534(.A1(new_n510_), .A2(new_n346_), .ZN(new_n721_));
  NAND2_X1  g535(.A1(new_n721_), .A2(new_n464_), .ZN(new_n722_));
  NAND2_X1  g536(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g537(.A(KEYINPUT83), .B1(new_n723_), .B2(new_n463_), .ZN(new_n724_));
  INV_X1    g538(.A(KEYINPUT83), .ZN(new_n725_));
  INV_X1    g539(.A(new_n463_), .ZN(new_n726_));
  AOI211_X1 g540(.A(new_n725_), .B(new_n726_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n727_));
  NOR2_X1   g541(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g542(.A1(new_n622_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g543(.A1(new_n717_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g544(.A(new_n730_), .B(new_n206_), .ZN(G15));
  NAND3_X1  g545(.A1(new_n641_), .A2(new_n350_), .A3(new_n667_), .ZN(new_n732_));
  NOR2_X1   g546(.A1(new_n732_), .A2(new_n729_), .ZN(new_n733_));
  INV_X1    g547(.A(KEYINPUT84), .ZN(new_n734_));
  XNOR2_X1  g548(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g549(.A(new_n735_), .B(G116), .ZN(G18));
  INV_X1    g550(.A(new_n728_), .ZN(new_n737_));
  INV_X1    g551(.A(new_n691_), .ZN(new_n738_));
  OR3_X1    g552(.A1(new_n462_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  XOR2_X1   g553(.A(KEYINPUT85), .B(G119), .Z(new_n740_));
  XNOR2_X1  g554(.A(new_n739_), .B(new_n740_), .ZN(G21));
  NOR2_X1   g555(.A1(new_n636_), .A2(new_n615_), .ZN(new_n742_));
  AND3_X1   g556(.A1(new_n728_), .A2(new_n742_), .A3(new_n704_), .ZN(new_n743_));
  AND3_X1   g557(.A1(new_n700_), .A2(KEYINPUT86), .A3(new_n351_), .ZN(new_n744_));
  AOI21_X1  g558(.A(KEYINPUT86), .B1(new_n700_), .B2(new_n351_), .ZN(new_n745_));
  OAI21_X1  g559(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g560(.A(new_n746_), .B(G122), .ZN(G24));
  NOR4_X1   g561(.A1(new_n679_), .A2(new_n423_), .A3(new_n658_), .A4(new_n687_), .ZN(new_n748_));
  NAND4_X1  g562(.A1(new_n331_), .A2(new_n728_), .A3(new_n748_), .A4(new_n336_), .ZN(new_n749_));
  XOR2_X1   g563(.A(KEYINPUT87), .B(G125), .Z(new_n750_));
  XNOR2_X1  g564(.A(new_n749_), .B(new_n750_), .ZN(G27));
  NOR2_X1   g565(.A1(new_n335_), .A2(new_n639_), .ZN(new_n752_));
  INV_X1    g566(.A(new_n752_), .ZN(new_n753_));
  NOR2_X1   g567(.A1(new_n753_), .A2(new_n523_), .ZN(new_n754_));
  NAND3_X1  g568(.A1(new_n754_), .A2(new_n622_), .A3(new_n714_), .ZN(new_n755_));
  XNOR2_X1  g569(.A(new_n755_), .B(G131), .ZN(G33));
  NAND3_X1  g570(.A1(new_n754_), .A2(new_n622_), .A3(new_n688_), .ZN(new_n757_));
  XNOR2_X1  g571(.A(new_n757_), .B(G134), .ZN(G36));
  OAI21_X1  g572(.A(new_n665_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n759_));
  NOR2_X1   g573(.A1(new_n759_), .A2(new_n690_), .ZN(new_n760_));
  INV_X1    g574(.A(new_n687_), .ZN(new_n761_));
  AOI21_X1  g575(.A(new_n502_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n762_));
  OAI211_X1 g576(.A(new_n505_), .B(new_n508_), .C1(KEYINPUT89), .C2(new_n762_), .ZN(new_n763_));
  AND2_X1   g577(.A1(new_n762_), .A2(KEYINPUT89), .ZN(new_n764_));
  AOI21_X1  g578(.A(KEYINPUT88), .B1(new_n507_), .B2(new_n492_), .ZN(new_n765_));
  NAND3_X1  g579(.A1(new_n507_), .A2(new_n492_), .A3(KEYINPUT88), .ZN(new_n766_));
  NAND2_X1  g580(.A1(new_n766_), .A2(new_n502_), .ZN(new_n767_));
  OAI22_X1  g581(.A1(new_n763_), .A2(new_n764_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g582(.A(new_n464_), .B1(new_n768_), .B2(new_n346_), .ZN(new_n769_));
  OAI211_X1 g583(.A(new_n463_), .B(new_n761_), .C1(new_n514_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g584(.A(new_n770_), .ZN(new_n771_));
  NAND4_X1  g585(.A1(new_n760_), .A2(new_n752_), .A3(new_n636_), .A4(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g586(.A(new_n772_), .B(G137), .ZN(G39));
  OAI21_X1  g587(.A(new_n463_), .B1(new_n514_), .B2(new_n769_), .ZN(new_n774_));
  XNOR2_X1  g588(.A(new_n774_), .B(KEYINPUT90), .ZN(new_n775_));
  NOR2_X1   g589(.A1(new_n619_), .A2(new_n620_), .ZN(new_n776_));
  NAND4_X1  g590(.A1(new_n775_), .A2(new_n714_), .A3(new_n752_), .A4(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g591(.A(new_n777_), .B(G140), .ZN(G42));
  AND4_X1   g592(.A1(new_n623_), .A2(new_n681_), .A3(new_n660_), .A4(new_n668_), .ZN(new_n779_));
  NAND2_X1  g593(.A1(new_n739_), .A2(new_n746_), .ZN(new_n780_));
  NOR2_X1   g594(.A1(new_n780_), .A2(new_n730_), .ZN(new_n781_));
  NAND3_X1  g595(.A1(new_n735_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g596(.A1(new_n715_), .A2(new_n749_), .ZN(new_n783_));
  XNOR2_X1  g597(.A(new_n783_), .B(KEYINPUT104), .ZN(new_n784_));
  NOR2_X1   g598(.A1(new_n523_), .A2(new_n687_), .ZN(new_n785_));
  NAND3_X1  g599(.A1(new_n641_), .A2(new_n711_), .A3(new_n785_), .ZN(new_n786_));
  AND2_X1   g600(.A1(new_n697_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g601(.A1(new_n784_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g602(.A1(new_n788_), .A2(KEYINPUT105), .ZN(new_n789_));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n790_));
  NAND3_X1  g604(.A1(new_n784_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g605(.A(new_n782_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g606(.A1(new_n755_), .A2(new_n757_), .ZN(new_n793_));
  INV_X1    g607(.A(KEYINPUT102), .ZN(new_n794_));
  NAND2_X1  g608(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g609(.A(new_n748_), .ZN(new_n796_));
  INV_X1    g610(.A(KEYINPUT100), .ZN(new_n797_));
  AOI21_X1  g611(.A(new_n796_), .B1(new_n754_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g612(.A(new_n798_), .B1(new_n797_), .B2(new_n754_), .ZN(new_n799_));
  XNOR2_X1  g613(.A(new_n460_), .B(KEYINPUT101), .ZN(new_n800_));
  NAND4_X1  g614(.A1(new_n785_), .A2(new_n800_), .A3(new_n691_), .A4(new_n752_), .ZN(new_n801_));
  NAND3_X1  g615(.A1(new_n795_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  NOR2_X1   g616(.A1(new_n793_), .A2(new_n794_), .ZN(new_n803_));
  OAI21_X1  g617(.A(KEYINPUT103), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AND2_X1   g618(.A1(new_n799_), .A2(new_n801_), .ZN(new_n805_));
  INV_X1    g619(.A(new_n803_), .ZN(new_n806_));
  INV_X1    g620(.A(KEYINPUT103), .ZN(new_n807_));
  NAND4_X1  g621(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .A4(new_n795_), .ZN(new_n808_));
  NAND2_X1  g622(.A1(new_n804_), .A2(new_n808_), .ZN(new_n809_));
  AND3_X1   g623(.A1(new_n792_), .A2(KEYINPUT106), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g624(.A(KEYINPUT106), .B1(new_n792_), .B2(new_n809_), .ZN(new_n811_));
  NOR2_X1   g625(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g626(.A1(new_n759_), .A2(new_n345_), .ZN(new_n813_));
  XNOR2_X1  g627(.A(new_n813_), .B(KEYINPUT93), .ZN(new_n814_));
  NAND2_X1  g628(.A1(new_n814_), .A2(new_n742_), .ZN(new_n815_));
  XNOR2_X1  g629(.A(new_n815_), .B(KEYINPUT96), .ZN(new_n816_));
  NOR4_X1   g630(.A1(new_n816_), .A2(new_n638_), .A3(new_n640_), .A4(new_n737_), .ZN(new_n817_));
  XNOR2_X1  g631(.A(new_n817_), .B(KEYINPUT97), .ZN(new_n818_));
  NAND3_X1  g632(.A1(new_n814_), .A2(new_n728_), .A3(new_n752_), .ZN(new_n819_));
  INV_X1    g633(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g634(.A1(new_n820_), .A2(new_n622_), .ZN(new_n821_));
  XNOR2_X1  g635(.A(new_n821_), .B(KEYINPUT94), .ZN(new_n822_));
  INV_X1    g636(.A(new_n423_), .ZN(new_n823_));
  NOR3_X1   g637(.A1(new_n335_), .A2(new_n823_), .A3(new_n710_), .ZN(new_n824_));
  XNOR2_X1  g638(.A(new_n824_), .B(KEYINPUT95), .ZN(new_n825_));
  NOR3_X1   g639(.A1(new_n658_), .A2(new_n615_), .A3(new_n639_), .ZN(new_n826_));
  NAND4_X1  g640(.A1(new_n825_), .A2(new_n463_), .A3(new_n723_), .A4(new_n826_), .ZN(new_n827_));
  NOR4_X1   g641(.A1(new_n753_), .A2(new_n615_), .A3(new_n345_), .A4(new_n710_), .ZN(new_n828_));
  NAND4_X1  g642(.A1(new_n828_), .A2(new_n423_), .A3(new_n658_), .A4(new_n728_), .ZN(new_n829_));
  XOR2_X1   g643(.A(new_n829_), .B(KEYINPUT99), .Z(new_n830_));
  NAND4_X1  g644(.A1(new_n822_), .A2(new_n340_), .A3(new_n827_), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g645(.A(KEYINPUT91), .ZN(new_n832_));
  NAND2_X1  g646(.A1(new_n659_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g647(.A(KEYINPUT91), .B1(new_n423_), .B2(new_n658_), .ZN(new_n834_));
  NAND2_X1  g648(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g649(.A1(new_n828_), .A2(new_n728_), .A3(new_n835_), .ZN(new_n836_));
  AOI22_X1  g650(.A1(new_n820_), .A2(new_n680_), .B1(new_n836_), .B2(KEYINPUT92), .ZN(new_n837_));
  AOI21_X1  g651(.A(new_n775_), .B1(new_n726_), .B2(new_n723_), .ZN(new_n838_));
  NOR2_X1   g652(.A1(new_n838_), .A2(new_n753_), .ZN(new_n839_));
  NOR2_X1   g653(.A1(new_n335_), .A2(new_n187_), .ZN(new_n840_));
  XOR2_X1   g654(.A(new_n840_), .B(KEYINPUT98), .Z(new_n841_));
  AOI21_X1  g655(.A(new_n839_), .B1(new_n728_), .B2(new_n841_), .ZN(new_n842_));
  OAI221_X1 g656(.A(new_n837_), .B1(KEYINPUT92), .B2(new_n836_), .C1(new_n816_), .C2(new_n842_), .ZN(new_n843_));
  NOR3_X1   g657(.A1(new_n818_), .A2(new_n831_), .A3(new_n843_), .ZN(new_n844_));
  NOR2_X1   g658(.A1(G952), .A2(G953), .ZN(new_n845_));
  AOI22_X1  g659(.A1(new_n812_), .A2(new_n844_), .B1(new_n827_), .B2(new_n845_), .ZN(G75));
  AOI211_X1 g660(.A(new_n309_), .B(new_n190_), .C1(new_n792_), .C2(new_n809_), .ZN(new_n847_));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n848_));
  XOR2_X1   g662(.A(new_n318_), .B(KEYINPUT108), .Z(new_n849_));
  XOR2_X1   g663(.A(new_n849_), .B(KEYINPUT107), .Z(new_n850_));
  XNOR2_X1  g664(.A(new_n850_), .B(new_n320_), .ZN(new_n851_));
  AND3_X1   g665(.A1(new_n847_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g666(.A(new_n851_), .B(new_n848_), .ZN(new_n853_));
  NOR2_X1   g667(.A1(new_n847_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g668(.A1(new_n339_), .A2(G952), .ZN(new_n855_));
  NOR3_X1   g669(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(G51));
  NAND2_X1  g670(.A1(G469), .A2(G902), .ZN(new_n857_));
  OAI22_X1  g671(.A1(new_n812_), .A2(new_n857_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n858_));
  NAND2_X1  g672(.A1(new_n792_), .A2(new_n809_), .ZN(new_n859_));
  OR2_X1    g673(.A1(new_n768_), .A2(new_n857_), .ZN(new_n860_));
  INV_X1    g674(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g675(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g676(.A(new_n855_), .B1(new_n858_), .B2(new_n862_), .ZN(G54));
  NAND3_X1  g677(.A1(new_n859_), .A2(G475), .A3(G902), .ZN(new_n864_));
  NAND2_X1  g678(.A1(new_n403_), .A2(new_n410_), .ZN(new_n865_));
  NAND2_X1  g679(.A1(new_n865_), .A2(KEYINPUT110), .ZN(new_n866_));
  NAND2_X1  g680(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g681(.A(new_n855_), .ZN(new_n868_));
  INV_X1    g682(.A(new_n866_), .ZN(new_n869_));
  NAND4_X1  g683(.A1(new_n859_), .A2(G475), .A3(G902), .A4(new_n869_), .ZN(new_n870_));
  NAND3_X1  g684(.A1(new_n867_), .A2(new_n868_), .A3(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g685(.A(new_n871_), .B(KEYINPUT111), .ZN(G60));
  MUX2_X1   g686(.A(new_n647_), .B(KEYINPUT69), .S(new_n648_), .Z(new_n873_));
  INV_X1    g687(.A(new_n812_), .ZN(new_n874_));
  NOR2_X1   g688(.A1(new_n424_), .A2(new_n346_), .ZN(new_n875_));
  AOI21_X1  g689(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g690(.A(new_n873_), .B(new_n875_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n877_));
  NAND2_X1  g691(.A1(new_n877_), .A2(new_n868_), .ZN(new_n878_));
  NOR2_X1   g692(.A1(new_n876_), .A2(new_n878_), .ZN(G63));
  NAND3_X1  g693(.A1(new_n859_), .A2(G217), .A3(new_n310_), .ZN(new_n880_));
  NOR3_X1   g694(.A1(new_n880_), .A2(KEYINPUT112), .A3(new_n672_), .ZN(new_n881_));
  AOI21_X1  g695(.A(new_n881_), .B1(new_n608_), .B2(new_n880_), .ZN(new_n882_));
  OAI21_X1  g696(.A(KEYINPUT112), .B1(new_n880_), .B2(new_n672_), .ZN(new_n883_));
  AOI21_X1  g697(.A(new_n855_), .B1(new_n882_), .B2(new_n883_), .ZN(G66));
  INV_X1    g698(.A(new_n782_), .ZN(new_n885_));
  OAI21_X1  g699(.A(KEYINPUT113), .B1(new_n885_), .B2(G953), .ZN(new_n886_));
  INV_X1    g700(.A(new_n339_), .ZN(new_n887_));
  AOI21_X1  g701(.A(new_n849_), .B1(new_n348_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g702(.A(KEYINPUT113), .ZN(new_n889_));
  NAND3_X1  g703(.A1(new_n782_), .A2(new_n889_), .A3(new_n282_), .ZN(new_n890_));
  NAND3_X1  g704(.A1(new_n886_), .A2(new_n888_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n892_));
  AND2_X1   g706(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g707(.A(new_n888_), .B1(new_n886_), .B2(new_n890_), .ZN(new_n894_));
  NOR2_X1   g708(.A1(new_n894_), .A2(KEYINPUT114), .ZN(new_n895_));
  NOR2_X1   g709(.A1(new_n891_), .A2(new_n892_), .ZN(new_n896_));
  NOR3_X1   g710(.A1(new_n893_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g711(.A(new_n282_), .B1(G224), .B2(G898), .ZN(new_n898_));
  AOI21_X1  g712(.A(new_n898_), .B1(new_n894_), .B2(KEYINPUT114), .ZN(new_n899_));
  AOI22_X1  g713(.A1(new_n897_), .A2(new_n899_), .B1(new_n898_), .B2(new_n888_), .ZN(G69));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n901_));
  XNOR2_X1  g715(.A(new_n544_), .B(KEYINPUT116), .ZN(new_n902_));
  NAND2_X1  g716(.A1(new_n902_), .A2(new_n377_), .ZN(new_n903_));
  NAND2_X1  g717(.A1(new_n684_), .A2(G953), .ZN(new_n904_));
  NAND2_X1  g718(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g719(.A1(new_n902_), .A2(new_n377_), .ZN(new_n906_));
  NOR2_X1   g720(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  AND2_X1   g721(.A1(new_n693_), .A2(new_n696_), .ZN(new_n908_));
  NAND2_X1  g722(.A1(new_n777_), .A2(new_n772_), .ZN(new_n909_));
  NOR4_X1   g723(.A1(new_n908_), .A2(new_n712_), .A3(new_n783_), .A4(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g724(.A(new_n666_), .B(KEYINPUT119), .ZN(new_n911_));
  NAND3_X1  g725(.A1(new_n911_), .A2(new_n834_), .A3(new_n833_), .ZN(new_n912_));
  AND2_X1   g726(.A1(new_n622_), .A2(new_n752_), .ZN(new_n913_));
  NAND3_X1  g727(.A1(new_n912_), .A2(new_n913_), .A3(new_n785_), .ZN(new_n914_));
  XOR2_X1   g728(.A(new_n914_), .B(KEYINPUT120), .Z(new_n915_));
  AOI211_X1 g729(.A(new_n887_), .B(new_n907_), .C1(new_n910_), .C2(new_n915_), .ZN(new_n916_));
  NAND4_X1  g730(.A1(new_n755_), .A2(new_n757_), .A3(new_n772_), .A4(new_n777_), .ZN(new_n917_));
  NOR3_X1   g731(.A1(new_n770_), .A2(new_n423_), .A3(new_n459_), .ZN(new_n918_));
  NAND4_X1  g732(.A1(new_n622_), .A2(new_n331_), .A3(new_n336_), .A4(new_n918_), .ZN(new_n919_));
  NAND3_X1  g733(.A1(new_n715_), .A2(new_n749_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g734(.A(new_n920_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n921_));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n922_));
  AOI21_X1  g736(.A(new_n917_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g737(.A(KEYINPUT117), .B1(new_n908_), .B2(new_n920_), .ZN(new_n924_));
  AOI21_X1  g738(.A(G953), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g739(.A(new_n907_), .ZN(new_n926_));
  OAI21_X1  g740(.A(KEYINPUT118), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  AND3_X1   g741(.A1(new_n715_), .A2(new_n749_), .A3(new_n919_), .ZN(new_n928_));
  NAND3_X1  g742(.A1(new_n697_), .A2(new_n928_), .A3(new_n922_), .ZN(new_n929_));
  NOR2_X1   g743(.A1(new_n793_), .A2(new_n909_), .ZN(new_n930_));
  NAND2_X1  g744(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  AOI21_X1  g745(.A(new_n922_), .B1(new_n697_), .B2(new_n928_), .ZN(new_n932_));
  OAI21_X1  g746(.A(new_n282_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g747(.A(KEYINPUT118), .ZN(new_n934_));
  NAND3_X1  g748(.A1(new_n933_), .A2(new_n934_), .A3(new_n907_), .ZN(new_n935_));
  AOI21_X1  g749(.A(new_n916_), .B1(new_n927_), .B2(new_n935_), .ZN(new_n936_));
  AOI21_X1  g750(.A(new_n339_), .B1(G227), .B2(G900), .ZN(new_n937_));
  OAI21_X1  g751(.A(new_n901_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g752(.A1(new_n910_), .A2(new_n915_), .ZN(new_n939_));
  NAND3_X1  g753(.A1(new_n939_), .A2(new_n339_), .A3(new_n926_), .ZN(new_n940_));
  NAND3_X1  g754(.A1(new_n924_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n941_));
  AOI211_X1 g755(.A(KEYINPUT118), .B(new_n926_), .C1(new_n941_), .C2(new_n282_), .ZN(new_n942_));
  AOI21_X1  g756(.A(new_n934_), .B1(new_n933_), .B2(new_n907_), .ZN(new_n943_));
  OAI21_X1  g757(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g758(.A(new_n937_), .ZN(new_n945_));
  NAND3_X1  g759(.A1(new_n944_), .A2(KEYINPUT121), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g760(.A1(new_n938_), .A2(new_n946_), .ZN(new_n947_));
  OAI211_X1 g761(.A(new_n937_), .B(new_n940_), .C1(new_n942_), .C2(new_n943_), .ZN(new_n948_));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949_));
  NAND2_X1  g763(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g764(.A1(new_n927_), .A2(new_n935_), .ZN(new_n951_));
  NAND4_X1  g765(.A1(new_n951_), .A2(KEYINPUT122), .A3(new_n937_), .A4(new_n940_), .ZN(new_n952_));
  NAND2_X1  g766(.A1(new_n950_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g767(.A1(new_n947_), .A2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g768(.A1(new_n954_), .A2(KEYINPUT123), .ZN(new_n955_));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n956_));
  NAND3_X1  g770(.A1(new_n947_), .A2(new_n953_), .A3(new_n956_), .ZN(new_n957_));
  NAND2_X1  g771(.A1(new_n955_), .A2(new_n957_), .ZN(G72));
  AOI21_X1  g772(.A(new_n585_), .B1(new_n792_), .B2(new_n809_), .ZN(new_n959_));
  NAND2_X1  g773(.A1(new_n565_), .A2(new_n566_), .ZN(new_n960_));
  XNOR2_X1  g774(.A(new_n960_), .B(KEYINPUT124), .ZN(new_n961_));
  OR3_X1    g775(.A1(new_n959_), .A2(KEYINPUT125), .A3(new_n961_), .ZN(new_n962_));
  OAI21_X1  g776(.A(KEYINPUT125), .B1(new_n959_), .B2(new_n961_), .ZN(new_n963_));
  OR2_X1    g777(.A1(new_n782_), .A2(new_n941_), .ZN(new_n964_));
  NAND2_X1  g778(.A1(new_n961_), .A2(new_n584_), .ZN(new_n965_));
  INV_X1    g779(.A(new_n965_), .ZN(new_n966_));
  AOI21_X1  g780(.A(new_n560_), .B1(new_n964_), .B2(new_n966_), .ZN(new_n967_));
  NAND3_X1  g781(.A1(new_n962_), .A2(new_n963_), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1  g782(.A(new_n965_), .B1(new_n792_), .B2(new_n809_), .ZN(new_n969_));
  NAND3_X1  g783(.A1(new_n910_), .A2(new_n915_), .A3(new_n779_), .ZN(new_n970_));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n971_));
  AOI21_X1  g785(.A(new_n971_), .B1(new_n735_), .B2(new_n781_), .ZN(new_n972_));
  NOR2_X1   g786(.A1(new_n970_), .A2(new_n972_), .ZN(new_n973_));
  NAND3_X1  g787(.A1(new_n735_), .A2(new_n781_), .A3(new_n971_), .ZN(new_n974_));
  AOI21_X1  g788(.A(new_n585_), .B1(new_n973_), .B2(new_n974_), .ZN(new_n975_));
  OAI22_X1  g789(.A1(new_n969_), .A2(KEYINPUT126), .B1(new_n975_), .B2(new_n961_), .ZN(new_n976_));
  AND2_X1   g790(.A1(new_n969_), .A2(KEYINPUT126), .ZN(new_n977_));
  OAI21_X1  g791(.A(new_n560_), .B1(new_n976_), .B2(new_n977_), .ZN(new_n978_));
  AND3_X1   g792(.A1(new_n968_), .A2(new_n978_), .A3(new_n868_), .ZN(G57));
endmodule


