//Secret key is'0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_c1355" written by ABC on Sun Nov 20 19:50:24 2022

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat,
    G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G134gat), .B(G162gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT32), .ZN(new_n208_));
  INV_X1    g007(.A(G43gat), .ZN(new_n209_));
  INV_X1    g008(.A(G50gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT33), .B(G43gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n210_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n207_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT34), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n208_), .A2(KEYINPUT34), .A3(new_n214_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT43), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(KEYINPUT43), .A3(new_n219_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n225_), .B(KEYINPUT19), .Z(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT17), .B1(G85gat), .B2(G92gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT22), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT22), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n229_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(new_n233_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT18), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n242_), .A2(new_n244_), .B1(G85gat), .B2(G92gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n225_), .B(KEYINPUT19), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n246_), .A2(KEYINPUT20), .B1(new_n227_), .B2(new_n228_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT20), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n226_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n245_), .A2(KEYINPUT21), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT21), .B1(new_n245_), .B2(new_n250_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n240_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT28), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n245_), .A2(new_n250_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n245_), .A2(new_n250_), .A3(KEYINPUT21), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n240_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n224_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n253_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n220_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(G232gat), .B(G233gat), .C1(new_n262_), .C2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n222_), .A2(new_n223_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n260_), .B1(new_n259_), .B2(new_n240_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n240_), .ZN(new_n270_));
  AOI211_X1 g069(.A(KEYINPUT28), .B(new_n270_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G232gat), .A2(G233gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n265_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n206_), .B1(new_n267_), .B2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n206_), .B(KEYINPUT85), .Z(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n272_), .B2(new_n265_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n274_), .B(new_n276_), .C1(new_n277_), .C2(KEYINPUT86), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n267_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT87), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n274_), .A2(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n267_), .A2(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(KEYINPUT86), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT87), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n275_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT64), .B(G183gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT65), .B1(new_n288_), .B2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290_));
  INV_X1    g089(.A(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(G183gat), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n292_), .A2(KEYINPUT64), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(KEYINPUT64), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n290_), .B(new_n291_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n292_), .A2(new_n291_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT63), .B1(G169gat), .B2(G176gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(KEYINPUT63), .A2(G169gat), .A3(G176gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(KEYINPUT62), .A2(G169gat), .A3(G176gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT62), .B1(G169gat), .B2(G176gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n297_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n296_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n296_), .A2(new_n305_), .A3(KEYINPUT66), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(KEYINPUT59), .A2(G176gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(KEYINPUT59), .A2(G176gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT60), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT60), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(new_n310_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n297_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT61), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT61), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n324_), .A3(new_n321_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n308_), .A2(new_n309_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(G113gat), .ZN(new_n327_));
  INV_X1    g126(.A(G120gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G113gat), .A2(G120gat), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G127gat), .A2(G134gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT3), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(G127gat), .A3(G134gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337_));
  INV_X1    g136(.A(G127gat), .ZN(new_n338_));
  INV_X1    g137(.A(G134gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n331_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n333_), .A2(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n337_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT12), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n337_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n344_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT2), .B1(new_n344_), .B2(new_n337_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n350_), .B(new_n351_), .C1(new_n352_), .C2(new_n331_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n326_), .A2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n347_), .A2(new_n353_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n296_), .A2(new_n305_), .A3(KEYINPUT66), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT66), .B1(new_n296_), .B2(new_n305_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n324_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n359_));
  AOI211_X1 g158(.A(KEYINPUT61), .B(new_n320_), .C1(new_n314_), .C2(new_n316_), .ZN(new_n360_));
  OAI22_X1  g159(.A1(new_n357_), .A2(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n355_), .A2(new_n362_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n355_), .A2(new_n362_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n364_), .B(new_n363_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT73), .Z(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n373_), .A2(KEYINPUT75), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n365_), .B(new_n371_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(KEYINPUT75), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT76), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n379_), .A3(new_n376_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT72), .ZN(new_n383_));
  AND3_X1   g182(.A1(KEYINPUT53), .A2(G197gat), .A3(G204gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT53), .B1(G197gat), .B2(G204gat), .ZN(new_n385_));
  OAI22_X1  g184(.A1(new_n384_), .A2(new_n385_), .B1(G197gat), .B2(G204gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT55), .ZN(new_n388_));
  INV_X1    g187(.A(G211gat), .ZN(new_n389_));
  INV_X1    g188(.A(G218gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT54), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT54), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G211gat), .A3(G218gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n386_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT57), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT56), .B(G218gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(new_n389_), .ZN(new_n399_));
  AND2_X1   g198(.A1(KEYINPUT56), .A2(G218gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT56), .A2(G218gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n397_), .B(new_n389_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n386_), .A2(new_n394_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT58), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n389_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT57), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n402_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT58), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n405_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n396_), .B1(new_n407_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n414_));
  INV_X1    g213(.A(G155gat), .ZN(new_n415_));
  INV_X1    g214(.A(G162gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT7), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT7), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(G155gat), .A3(G162gat), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n417_), .A2(KEYINPUT8), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT8), .B1(new_n417_), .B2(new_n419_), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n420_), .A2(new_n421_), .B1(G155gat), .B2(G162gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT6), .B(G141gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n422_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT11), .ZN(new_n430_));
  OR2_X1    g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n417_), .A2(new_n419_), .B1(new_n431_), .B2(new_n423_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT9), .B(G155gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n416_), .ZN(new_n435_));
  AND2_X1   g234(.A1(KEYINPUT9), .A2(G155gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(KEYINPUT9), .A2(G155gat), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n433_), .B(new_n416_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n430_), .B(new_n432_), .C1(new_n435_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n416_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT10), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n438_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n430_), .B1(new_n444_), .B2(new_n432_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n414_), .B(new_n429_), .C1(new_n441_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n432_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT11), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n440_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n414_), .B1(new_n450_), .B2(new_n429_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n413_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n429_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT71), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n404_), .A2(KEYINPUT58), .A3(new_n406_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n411_), .B1(new_n410_), .B2(new_n405_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n395_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n459_), .A3(new_n446_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n452_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT70), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n454_), .B1(new_n452_), .B2(new_n460_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n383_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n452_), .A2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n453_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n383_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(KEYINPUT70), .A3(new_n467_), .A4(new_n461_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G78gat), .B(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n470_), .A3(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(new_n235_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT0), .B(G57gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n449_), .A2(new_n440_), .B1(new_n422_), .B2(new_n428_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n356_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n354_), .A2(new_n455_), .A3(KEYINPUT13), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n350_), .B1(new_n352_), .B2(new_n331_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(new_n429_), .C1(new_n441_), .C2(new_n445_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n450_), .A2(KEYINPUT14), .A3(new_n429_), .A4(new_n487_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n486_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(KEYINPUT15), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n487_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n455_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n488_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n485_), .B(KEYINPUT1), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT15), .B1(new_n484_), .B2(new_n492_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n479_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n484_), .A2(new_n492_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n505_), .A2(new_n478_), .A3(new_n499_), .A4(new_n493_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n361_), .B2(new_n413_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n308_), .A2(new_n309_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n323_), .A2(new_n325_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n459_), .A2(new_n510_), .A3(KEYINPUT67), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n361_), .A2(new_n413_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G226gat), .A2(G233gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT52), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT68), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n515_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n361_), .A2(new_n413_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(new_n513_), .A3(KEYINPUT68), .A4(new_n515_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT50), .B(KEYINPUT51), .Z(new_n525_));
  XNOR2_X1  g324(.A(G64gat), .B(G92gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G8gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n517_), .A2(new_n521_), .A3(new_n523_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(KEYINPUT69), .A3(new_n532_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n507_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n381_), .A2(KEYINPUT77), .A3(new_n474_), .A4(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT77), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n378_), .A2(new_n474_), .A3(new_n380_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT78), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n532_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n530_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n524_), .A2(new_n545_), .A3(new_n529_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n507_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT79), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n482_), .A2(new_n483_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n490_), .A2(new_n491_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n550_), .B(new_n486_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n482_), .A2(new_n483_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT79), .B1(new_n554_), .B2(new_n485_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n495_), .A2(new_n488_), .A3(new_n497_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT80), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n479_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n533_), .A3(new_n506_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n549_), .A2(new_n560_), .B1(new_n473_), .B2(new_n472_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT81), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n472_), .A2(new_n473_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n561_), .A2(new_n562_), .B1(new_n563_), .B2(new_n537_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n549_), .A2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n474_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT81), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n381_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT82), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT82), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n571_), .B(new_n381_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n544_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G57gat), .ZN(new_n574_));
  INV_X1    g373(.A(G64gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT26), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT26), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n577_), .B(new_n578_), .C1(G57gat), .C2(G64gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT23), .Z(new_n581_));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n581_), .A2(KEYINPUT24), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n580_), .B(KEYINPUT23), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT24), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n582_), .B(KEYINPUT25), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G57gat), .B(G64gat), .Z(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n584_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT39), .B(G22gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT38), .B(G15gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G1gat), .A2(G8gat), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(KEYINPUT37), .A2(G1gat), .A3(G8gat), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n600_), .C1(G1gat), .C2(G8gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G15gat), .A2(G22gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT40), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n596_), .A2(new_n605_), .A3(new_n601_), .A4(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(G15gat), .A2(G22gat), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n602_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n609_), .B2(new_n602_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT35), .B(G1gat), .ZN(new_n612_));
  INV_X1    g411(.A(G8gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n597_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n607_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n593_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT48), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT47), .Z(new_n620_));
  INV_X1    g419(.A(new_n593_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n615_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT44), .ZN(new_n624_));
  OAI221_X1 g423(.A(new_n618_), .B1(KEYINPUT49), .B2(new_n620_), .C1(new_n621_), .C2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G183gat), .B(G211gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT45), .B(KEYINPUT46), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n625_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n620_), .A2(KEYINPUT49), .ZN(new_n630_));
  XOR2_X1   g429(.A(G127gat), .B(G155gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n632_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636_));
  INV_X1    g435(.A(G204gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT16), .B(G176gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n638_), .B(new_n639_), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n263_), .A2(new_n621_), .ZN(new_n641_));
  INV_X1    g440(.A(G230gat), .ZN(new_n642_));
  INV_X1    g441(.A(G233gat), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n641_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n593_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT29), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n254_), .A2(new_n261_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT29), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n593_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n646_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n253_), .A2(new_n593_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT27), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n645_), .B1(new_n654_), .B2(new_n641_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n640_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n646_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n650_), .B1(new_n649_), .B2(new_n593_), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT29), .B(new_n621_), .C1(new_n254_), .C2(new_n261_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT27), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n653_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n641_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n644_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n640_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n656_), .A2(KEYINPUT30), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT30), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n640_), .C1(new_n652_), .C2(new_n655_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(G113gat), .B(G141gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(G169gat), .B(G197gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT31), .Z(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n616_), .B2(new_n220_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n616_), .A2(new_n220_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n264_), .B2(new_n623_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n616_), .A2(new_n220_), .A3(KEYINPUT41), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n677_), .A2(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(G229gat), .A2(G233gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n624_), .A2(new_n224_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n685_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n678_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n676_), .B1(new_n686_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n616_), .B(KEYINPUT44), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n678_), .B1(new_n691_), .B2(new_n268_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n685_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n693_), .B(new_n675_), .C1(new_n685_), .C2(new_n684_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n671_), .A2(new_n696_), .ZN(new_n697_));
  AND4_X1   g496(.A1(new_n287_), .A2(new_n573_), .A3(new_n635_), .A4(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n507_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G1gat), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT89), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n573_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n565_), .A2(new_n562_), .A3(new_n474_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n563_), .A2(new_n537_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n561_), .A2(new_n562_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n569_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n571_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n568_), .A2(KEYINPUT82), .A3(new_n569_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n543_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT89), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n696_), .B1(new_n703_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT90), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n281_), .A2(new_n286_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n275_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT90), .B(new_n275_), .C1(new_n281_), .C2(new_n286_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n713_), .A2(new_n635_), .A3(new_n670_), .A4(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n507_), .B(KEYINPUT88), .Z(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n612_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n701_), .B1(new_n721_), .B2(new_n724_), .ZN(G1324gat));
  NAND2_X1  g524(.A1(new_n535_), .A2(new_n536_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G8gat), .B1(new_n699_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n726_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n613_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n721_), .B2(new_n729_), .ZN(G1325gat));
  NAND2_X1  g529(.A1(new_n381_), .A2(new_n595_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n721_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT91), .ZN(new_n733_));
  OAI21_X1  g532(.A(G15gat), .B1(new_n699_), .B2(new_n569_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1326gat));
  NAND2_X1  g534(.A1(new_n563_), .A2(new_n594_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n721_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT93), .ZN(new_n738_));
  OAI21_X1  g537(.A(G22gat), .B1(new_n699_), .B2(new_n474_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT92), .Z(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1327gat));
  INV_X1    g540(.A(G29gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT94), .B1(new_n711_), .B2(new_n720_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT94), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n573_), .A2(new_n744_), .A3(new_n719_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n635_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n697_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n747_), .B2(new_n507_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n635_), .A2(new_n671_), .A3(new_n287_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n713_), .A2(new_n749_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n750_), .A2(G29gat), .A3(new_n722_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1328gat));
  INV_X1    g551(.A(G36gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n747_), .B2(new_n728_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n750_), .A2(G36gat), .A3(new_n726_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1329gat));
  NAND3_X1  g555(.A1(new_n746_), .A2(new_n381_), .A3(new_n697_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT95), .A3(G43gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT95), .B1(new_n757_), .B2(G43gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n381_), .A2(new_n212_), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n758_), .A2(new_n759_), .B1(new_n750_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT96), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1330gat));
  NOR3_X1   g562(.A1(new_n750_), .A2(G50gat), .A3(new_n474_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n747_), .A2(new_n563_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(G50gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT97), .ZN(G1331gat));
  AND2_X1   g566(.A1(new_n671_), .A2(KEYINPUT98), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n671_), .A2(KEYINPUT98), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n695_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n772_));
  AND4_X1   g571(.A1(new_n287_), .A2(new_n573_), .A3(new_n771_), .A4(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n507_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G57gat), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT99), .Z(new_n776_));
  INV_X1    g575(.A(KEYINPUT101), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n703_), .A2(new_n712_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n720_), .A3(new_n772_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT100), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n771_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n723_), .A2(new_n574_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n776_), .B(new_n777_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n779_), .B(KEYINPUT100), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n770_), .A3(new_n783_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n775_), .B(KEYINPUT99), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT101), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(G1332gat));
  NOR2_X1   g588(.A1(new_n770_), .A2(new_n726_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n575_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n773_), .A2(new_n728_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n785_), .A2(new_n791_), .B1(new_n575_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT102), .ZN(G1333gat));
  INV_X1    g593(.A(G71gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n773_), .B2(new_n381_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT103), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n381_), .A2(new_n795_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n782_), .B2(new_n798_), .ZN(G1334gat));
  INV_X1    g598(.A(G78gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n773_), .B2(new_n563_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT104), .Z(new_n802_));
  NAND2_X1  g601(.A1(new_n563_), .A2(new_n800_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n782_), .B2(new_n803_), .ZN(G1335gat));
  INV_X1    g603(.A(new_n635_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n287_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n696_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n709_), .A2(new_n710_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT89), .B1(new_n809_), .B2(new_n544_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n702_), .B(new_n543_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT105), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT105), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n778_), .A2(new_n814_), .A3(new_n808_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n770_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n235_), .A3(new_n723_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n770_), .A2(new_n695_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n746_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G85gat), .B1(new_n819_), .B2(new_n700_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT106), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1336gat));
  NAND2_X1  g622(.A1(new_n813_), .A2(new_n815_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n236_), .A3(new_n790_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G92gat), .B1(new_n819_), .B2(new_n726_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1337gat));
  NOR3_X1   g626(.A1(new_n819_), .A2(new_n227_), .A3(new_n569_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n816_), .A2(new_n381_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n227_), .ZN(G1338gat));
  NAND2_X1  g629(.A1(new_n743_), .A2(new_n745_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(new_n563_), .A3(new_n805_), .A4(new_n818_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G106gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT107), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT107), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n835_), .A3(G106gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n474_), .A2(G106gat), .ZN(new_n838_));
  AND4_X1   g637(.A1(KEYINPUT108), .A2(new_n824_), .A3(new_n771_), .A4(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT108), .B1(new_n816_), .B2(new_n838_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT109), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n837_), .B(new_n843_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1339gat));
  NOR2_X1   g644(.A1(new_n722_), .A2(new_n728_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n694_), .A2(new_n848_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n684_), .A2(new_n685_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT111), .A3(new_n693_), .A4(new_n675_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT112), .B1(new_n692_), .B2(new_n685_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n688_), .C1(new_n687_), .C2(new_n678_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n684_), .A2(new_n685_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n849_), .A2(new_n851_), .B1(new_n674_), .B2(new_n856_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n667_), .A2(new_n857_), .A3(new_n669_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n695_), .A2(new_n666_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n652_), .A2(KEYINPUT110), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n660_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n663_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n860_), .B(new_n862_), .C1(new_n645_), .C2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n859_), .B1(new_n864_), .B2(new_n640_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n287_), .B1(new_n858_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n857_), .A2(new_n666_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n640_), .B2(new_n864_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(KEYINPUT113), .A2(new_n866_), .B1(new_n719_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n287_), .C1(new_n858_), .C2(new_n865_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n635_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n772_), .B(new_n670_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n474_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n875_), .A2(KEYINPUT114), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(KEYINPUT114), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n569_), .B(new_n847_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G113gat), .B1(new_n879_), .B2(new_n696_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n866_), .A2(KEYINPUT113), .ZN(new_n883_));
  INV_X1    g682(.A(new_n717_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n718_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n868_), .A3(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n871_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n805_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(KEYINPUT115), .A3(new_n873_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n882_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n540_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n846_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n327_), .A3(new_n695_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n880_), .A2(new_n895_), .ZN(G1340gat));
  AOI21_X1  g695(.A(new_n328_), .B1(new_n878_), .B2(new_n671_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT116), .B(G120gat), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n893_), .A2(new_n770_), .A3(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n898_), .A2(new_n900_), .A3(KEYINPUT117), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n893_), .A2(new_n770_), .A3(new_n899_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n897_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1341gat));
  OAI21_X1  g704(.A(G127gat), .B1(new_n879_), .B2(new_n805_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n894_), .A2(new_n338_), .A3(new_n635_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1342gat));
  NAND3_X1  g707(.A1(new_n894_), .A2(new_n339_), .A3(new_n806_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n878_), .A2(new_n719_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(G134gat), .ZN(new_n912_));
  AOI211_X1 g711(.A(KEYINPUT118), .B(new_n339_), .C1(new_n878_), .C2(new_n719_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n909_), .B1(new_n912_), .B2(new_n913_), .ZN(G1343gat));
  NOR2_X1   g713(.A1(new_n381_), .A2(new_n474_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n888_), .B2(new_n873_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n846_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G141gat), .B1(new_n918_), .B2(new_n696_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT119), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n890_), .A2(new_n846_), .A3(new_n915_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n695_), .A2(new_n427_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1344gat));
  OAI21_X1  g722(.A(G148gat), .B1(new_n918_), .B2(new_n670_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n771_), .A2(new_n426_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n921_), .B2(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT120), .ZN(G1345gat));
  OAI21_X1  g726(.A(G155gat), .B1(new_n918_), .B2(new_n805_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n635_), .A2(new_n434_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n921_), .B2(new_n929_), .ZN(G1346gat));
  NOR3_X1   g729(.A1(new_n921_), .A2(G162gat), .A3(new_n287_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT121), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n917_), .A2(new_n719_), .A3(new_n846_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(G162gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n932_), .B1(new_n931_), .B2(new_n935_), .ZN(G1347gat));
  NAND2_X1  g735(.A1(new_n892_), .A2(new_n700_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n726_), .A2(new_n696_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n310_), .ZN(new_n939_));
  OR3_X1    g738(.A1(new_n937_), .A2(KEYINPUT122), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n876_), .A2(new_n877_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n726_), .A2(new_n507_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n941_), .A2(new_n381_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G169gat), .B1(new_n943_), .B2(new_n696_), .ZN(new_n944_));
  OAI21_X1  g743(.A(KEYINPUT122), .B1(new_n937_), .B2(new_n939_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n940_), .A2(new_n944_), .A3(new_n945_), .ZN(G1348gat));
  OAI21_X1  g745(.A(G176gat), .B1(new_n943_), .B2(new_n670_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n790_), .B1(new_n312_), .B2(new_n311_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n937_), .B2(new_n948_), .ZN(G1349gat));
  OAI21_X1  g748(.A(G183gat), .B1(new_n943_), .B2(new_n805_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n635_), .A2(new_n728_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n951_), .A2(new_n288_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n950_), .B1(new_n937_), .B2(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n943_), .B2(new_n720_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n287_), .A2(new_n726_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n291_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n937_), .B2(new_n956_), .ZN(G1351gat));
  AOI21_X1  g756(.A(KEYINPUT115), .B1(new_n888_), .B2(new_n873_), .ZN(new_n958_));
  AOI211_X1 g757(.A(new_n881_), .B(new_n874_), .C1(new_n887_), .C2(new_n805_), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n700_), .B(new_n915_), .C1(new_n958_), .C2(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n890_), .A2(KEYINPUT123), .A3(new_n700_), .A4(new_n915_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(G197gat), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n964_), .A2(new_n965_), .A3(new_n938_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n917_), .A2(new_n942_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967_), .B2(new_n696_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1352gat));
  OAI21_X1  g768(.A(G204gat), .B1(new_n967_), .B2(new_n670_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n970_), .B(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n790_), .A2(new_n637_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n973_), .ZN(new_n974_));
  AOI21_X1  g773(.A(KEYINPUT125), .B1(new_n964_), .B2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976_));
  AOI211_X1 g775(.A(new_n976_), .B(new_n973_), .C1(new_n962_), .C2(new_n963_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n972_), .B1(new_n975_), .B2(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  OAI211_X1 g779(.A(KEYINPUT126), .B(new_n972_), .C1(new_n975_), .C2(new_n977_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1353gat));
  NOR2_X1   g781(.A1(new_n951_), .A2(G211gat), .ZN(new_n983_));
  AND2_X1   g782(.A1(new_n964_), .A2(new_n983_), .ZN(new_n984_));
  OR2_X1    g783(.A1(new_n984_), .A2(KEYINPUT127), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(KEYINPUT127), .ZN(new_n986_));
  OAI21_X1  g785(.A(G211gat), .B1(new_n967_), .B2(new_n805_), .ZN(new_n987_));
  NAND3_X1  g786(.A1(new_n985_), .A2(new_n986_), .A3(new_n987_), .ZN(G1354gat));
  NAND3_X1  g787(.A1(new_n964_), .A2(new_n398_), .A3(new_n955_), .ZN(new_n989_));
  OAI21_X1  g788(.A(G218gat), .B1(new_n967_), .B2(new_n720_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n989_), .A2(new_n990_), .ZN(G1355gat));
endmodule


