//Secret key is'0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_c3540" written by ABC on Wed Oct 26 14:05:58 2022

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41,
    G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132,
    G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226,
    G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311,
    G317, G322, G326, G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13,
    G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124,
    G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213,
    G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283,
    G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137_, new_n138_, new_n139_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_;
  INV_X1    g000(.A(G58), .ZN(new_n137_));
  INV_X1    g001(.A(G68), .ZN(new_n138_));
  NAND2_X1  g002(.A1(new_n137_), .A2(new_n138_), .ZN(new_n139_));
  NOR3_X1   g003(.A1(new_n139_), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g005(.A1(G1), .A2(G20), .ZN(new_n142_));
  NOR2_X1   g006(.A1(new_n142_), .A2(G13), .ZN(new_n143_));
  INV_X1    g007(.A(new_n143_), .ZN(new_n144_));
  OAI21_X1  g008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n145_));
  NAND2_X1  g009(.A1(new_n139_), .A2(G50), .ZN(new_n146_));
  NAND3_X1  g010(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n147_));
  OAI22_X1  g011(.A1(new_n144_), .A2(new_n145_), .B1(new_n146_), .B2(new_n147_), .ZN(new_n148_));
  AOI22_X1  g012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n149_));
  AOI22_X1  g013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n150_));
  AOI22_X1  g014(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n151_));
  AOI22_X1  g015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n152_));
  NAND4_X1  g016(.A1(new_n149_), .A2(new_n150_), .A3(new_n151_), .A4(new_n152_), .ZN(new_n153_));
  AOI21_X1  g017(.A(new_n148_), .B1(new_n142_), .B2(new_n153_), .ZN(G361));
  XNOR2_X1  g018(.A(G264), .B(G270), .ZN(new_n155_));
  XNOR2_X1  g019(.A(new_n155_), .B(KEYINPUT0), .ZN(new_n156_));
  XNOR2_X1  g020(.A(G250), .B(G257), .ZN(new_n157_));
  XNOR2_X1  g021(.A(new_n156_), .B(new_n157_), .ZN(new_n158_));
  XOR2_X1   g022(.A(G226), .B(G232), .Z(new_n159_));
  XNOR2_X1  g023(.A(G238), .B(G244), .ZN(new_n160_));
  XNOR2_X1  g024(.A(new_n159_), .B(new_n160_), .ZN(new_n161_));
  XNOR2_X1  g025(.A(new_n158_), .B(new_n161_), .ZN(G358));
  XNOR2_X1  g026(.A(G68), .B(G77), .ZN(new_n163_));
  XNOR2_X1  g027(.A(G50), .B(G58), .ZN(new_n164_));
  XNOR2_X1  g028(.A(new_n163_), .B(new_n164_), .ZN(new_n165_));
  XOR2_X1   g029(.A(new_n165_), .B(KEYINPUT2), .Z(new_n166_));
  XNOR2_X1  g030(.A(G87), .B(G97), .ZN(new_n167_));
  INV_X1    g031(.A(G107), .ZN(new_n168_));
  XNOR2_X1  g032(.A(new_n167_), .B(new_n168_), .ZN(new_n169_));
  XOR2_X1   g033(.A(KEYINPUT1), .B(G116), .Z(new_n170_));
  XNOR2_X1  g034(.A(new_n169_), .B(new_n170_), .ZN(new_n171_));
  XNOR2_X1  g035(.A(new_n166_), .B(new_n171_), .ZN(G351));
  INV_X1    g036(.A(G41), .ZN(new_n173_));
  INV_X1    g037(.A(G45), .ZN(new_n174_));
  AOI21_X1  g038(.A(G1), .B1(new_n173_), .B2(new_n174_), .ZN(new_n175_));
  INV_X1    g039(.A(new_n175_), .ZN(new_n176_));
  AND2_X1   g040(.A1(G33), .A2(G41), .ZN(new_n177_));
  NAND2_X1  g041(.A1(G1), .A2(G13), .ZN(new_n178_));
  OAI21_X1  g042(.A(G274), .B1(new_n177_), .B2(new_n178_), .ZN(new_n179_));
  NOR2_X1   g043(.A1(new_n176_), .A2(new_n179_), .ZN(new_n180_));
  NOR2_X1   g044(.A1(new_n177_), .A2(new_n178_), .ZN(new_n181_));
  NOR2_X1   g045(.A1(new_n181_), .A2(new_n175_), .ZN(new_n182_));
  AOI21_X1  g046(.A(new_n180_), .B1(G226), .B2(new_n182_), .ZN(new_n183_));
  NOR2_X1   g047(.A1(G33), .A2(G1698), .ZN(new_n184_));
  NAND2_X1  g048(.A1(new_n184_), .A2(G222), .ZN(new_n185_));
  NAND2_X1  g049(.A1(G33), .A2(G77), .ZN(new_n186_));
  INV_X1    g050(.A(G223), .ZN(new_n187_));
  INV_X1    g051(.A(G33), .ZN(new_n188_));
  NAND2_X1  g052(.A1(new_n188_), .A2(G1698), .ZN(new_n189_));
  OAI211_X1 g053(.A(new_n185_), .B(new_n186_), .C1(new_n187_), .C2(new_n189_), .ZN(new_n190_));
  NAND2_X1  g054(.A1(new_n190_), .A2(new_n181_), .ZN(new_n191_));
  NAND2_X1  g055(.A1(new_n183_), .A2(new_n191_), .ZN(new_n192_));
  INV_X1    g056(.A(G169), .ZN(new_n193_));
  NAND2_X1  g057(.A1(new_n192_), .A2(new_n193_), .ZN(new_n194_));
  OAI21_X1  g058(.A(G20), .B1(new_n139_), .B2(G50), .ZN(new_n195_));
  NOR2_X1   g059(.A1(G20), .A2(G33), .ZN(new_n196_));
  NAND2_X1  g060(.A1(new_n196_), .A2(G150), .ZN(new_n197_));
  INV_X1    g061(.A(G20), .ZN(new_n198_));
  NAND2_X1  g062(.A1(new_n198_), .A2(G33), .ZN(new_n199_));
  OAI211_X1 g063(.A(new_n195_), .B(new_n197_), .C1(new_n137_), .C2(new_n199_), .ZN(new_n200_));
  NAND3_X1  g064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n201_));
  NAND2_X1  g065(.A1(new_n201_), .A2(new_n178_), .ZN(new_n202_));
  INV_X1    g066(.A(G50), .ZN(new_n203_));
  INV_X1    g067(.A(G1), .ZN(new_n204_));
  NAND3_X1  g068(.A1(new_n204_), .A2(G13), .A3(G20), .ZN(new_n205_));
  INV_X1    g069(.A(new_n205_), .ZN(new_n206_));
  AOI22_X1  g070(.A1(new_n200_), .A2(new_n202_), .B1(new_n203_), .B2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g071(.A1(new_n205_), .A2(new_n178_), .A3(new_n201_), .ZN(new_n208_));
  INV_X1    g072(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g073(.A1(new_n204_), .A2(G20), .ZN(new_n210_));
  NAND3_X1  g074(.A1(new_n209_), .A2(G50), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g075(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g076(.A(new_n194_), .B(new_n212_), .C1(G179), .C2(new_n192_), .ZN(new_n213_));
  NAND2_X1  g077(.A1(new_n192_), .A2(G200), .ZN(new_n214_));
  AND2_X1   g078(.A1(new_n207_), .A2(new_n211_), .ZN(new_n215_));
  NAND2_X1  g079(.A1(new_n182_), .A2(G226), .ZN(new_n216_));
  OAI211_X1 g080(.A(G1), .B(G13), .C1(new_n188_), .C2(new_n173_), .ZN(new_n217_));
  NAND3_X1  g081(.A1(new_n217_), .A2(G274), .A3(new_n175_), .ZN(new_n218_));
  NAND4_X1  g082(.A1(new_n216_), .A2(new_n191_), .A3(G190), .A4(new_n218_), .ZN(new_n219_));
  NAND4_X1  g083(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT9), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g084(.A(KEYINPUT9), .ZN(new_n221_));
  NAND3_X1  g085(.A1(new_n219_), .A2(new_n207_), .A3(new_n211_), .ZN(new_n222_));
  INV_X1    g086(.A(G200), .ZN(new_n223_));
  AOI21_X1  g087(.A(new_n223_), .B1(new_n183_), .B2(new_n191_), .ZN(new_n224_));
  OAI21_X1  g088(.A(new_n221_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g089(.A1(new_n213_), .A2(new_n220_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g090(.A(KEYINPUT12), .ZN(new_n227_));
  NAND2_X1  g091(.A1(G33), .A2(G87), .ZN(new_n228_));
  INV_X1    g092(.A(G226), .ZN(new_n229_));
  INV_X1    g093(.A(G1698), .ZN(new_n230_));
  NAND2_X1  g094(.A1(new_n188_), .A2(new_n230_), .ZN(new_n231_));
  OAI221_X1 g095(.A(new_n228_), .B1(new_n189_), .B2(new_n229_), .C1(new_n187_), .C2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g096(.A1(new_n232_), .A2(new_n181_), .ZN(new_n233_));
  NAND2_X1  g097(.A1(new_n182_), .A2(G232), .ZN(new_n234_));
  NAND3_X1  g098(.A1(new_n233_), .A2(new_n218_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g099(.A(G190), .ZN(new_n236_));
  OAI21_X1  g100(.A(new_n227_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g101(.A(new_n180_), .B1(G232), .B2(new_n182_), .ZN(new_n238_));
  NAND4_X1  g102(.A1(new_n238_), .A2(KEYINPUT12), .A3(G190), .A4(new_n233_), .ZN(new_n239_));
  NAND2_X1  g103(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g104(.A1(new_n209_), .A2(G58), .A3(new_n210_), .ZN(new_n241_));
  NAND2_X1  g105(.A1(new_n196_), .A2(G159), .ZN(new_n242_));
  OAI21_X1  g106(.A(new_n242_), .B1(new_n138_), .B2(new_n199_), .ZN(new_n243_));
  NAND2_X1  g107(.A1(G58), .A2(G68), .ZN(new_n244_));
  AOI21_X1  g108(.A(new_n198_), .B1(new_n139_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g109(.A(new_n202_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g110(.A1(new_n206_), .A2(new_n137_), .ZN(new_n247_));
  NAND3_X1  g111(.A1(new_n241_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g112(.A(new_n248_), .B1(new_n235_), .B2(G200), .ZN(new_n249_));
  AND2_X1   g113(.A1(new_n246_), .A2(new_n247_), .ZN(new_n250_));
  AOI22_X1  g114(.A1(new_n193_), .A2(new_n235_), .B1(new_n250_), .B2(new_n241_), .ZN(new_n251_));
  INV_X1    g115(.A(G179), .ZN(new_n252_));
  NAND3_X1  g116(.A1(new_n238_), .A2(new_n252_), .A3(new_n233_), .ZN(new_n253_));
  AOI22_X1  g117(.A1(new_n240_), .A2(new_n249_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g118(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g119(.A1(new_n182_), .A2(G244), .ZN(new_n256_));
  NAND2_X1  g120(.A1(new_n256_), .A2(KEYINPUT11), .ZN(new_n257_));
  INV_X1    g121(.A(KEYINPUT11), .ZN(new_n258_));
  NAND3_X1  g122(.A1(new_n182_), .A2(new_n258_), .A3(G244), .ZN(new_n259_));
  NAND2_X1  g123(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g124(.A1(G33), .A2(G107), .ZN(new_n261_));
  INV_X1    g125(.A(G238), .ZN(new_n262_));
  INV_X1    g126(.A(G232), .ZN(new_n263_));
  OAI221_X1 g127(.A(new_n261_), .B1(new_n189_), .B2(new_n262_), .C1(new_n263_), .C2(new_n231_), .ZN(new_n264_));
  AOI21_X1  g128(.A(new_n180_), .B1(new_n264_), .B2(new_n181_), .ZN(new_n265_));
  NAND2_X1  g129(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g130(.A1(new_n266_), .A2(G200), .ZN(new_n267_));
  OR2_X1    g131(.A1(new_n208_), .A2(KEYINPUT10), .ZN(new_n268_));
  NAND2_X1  g132(.A1(new_n208_), .A2(KEYINPUT10), .ZN(new_n269_));
  NAND4_X1  g133(.A1(new_n268_), .A2(G77), .A3(new_n210_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g134(.A(new_n202_), .ZN(new_n271_));
  NOR2_X1   g135(.A1(new_n198_), .A2(G77), .ZN(new_n272_));
  NOR2_X1   g136(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g137(.A(new_n228_), .B(new_n198_), .C1(G33), .C2(new_n137_), .ZN(new_n274_));
  INV_X1    g138(.A(G13), .ZN(new_n275_));
  NOR2_X1   g139(.A1(new_n275_), .A2(G1), .ZN(new_n276_));
  AOI22_X1  g140(.A1(new_n273_), .A2(new_n274_), .B1(new_n276_), .B2(new_n272_), .ZN(new_n277_));
  NAND3_X1  g141(.A1(new_n260_), .A2(G190), .A3(new_n265_), .ZN(new_n278_));
  NAND4_X1  g142(.A1(new_n267_), .A2(new_n270_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g143(.A1(new_n266_), .A2(new_n193_), .ZN(new_n280_));
  NAND2_X1  g144(.A1(new_n270_), .A2(new_n277_), .ZN(new_n281_));
  NAND3_X1  g145(.A1(new_n260_), .A2(new_n252_), .A3(new_n265_), .ZN(new_n282_));
  NAND3_X1  g146(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g147(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g148(.A1(new_n182_), .A2(G238), .ZN(new_n285_));
  INV_X1    g149(.A(G97), .ZN(new_n286_));
  OAI22_X1  g150(.A1(new_n189_), .A2(new_n263_), .B1(new_n188_), .B2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g151(.A1(new_n231_), .A2(new_n229_), .ZN(new_n288_));
  OAI21_X1  g152(.A(new_n181_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g153(.A1(new_n285_), .A2(new_n218_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g154(.A1(new_n290_), .A2(G200), .ZN(new_n291_));
  NAND4_X1  g155(.A1(new_n268_), .A2(G68), .A3(new_n210_), .A4(new_n269_), .ZN(new_n292_));
  AOI211_X1 g156(.A(new_n198_), .B(G68), .C1(new_n201_), .C2(new_n275_), .ZN(new_n293_));
  NAND2_X1  g157(.A1(new_n188_), .A2(G50), .ZN(new_n294_));
  AOI21_X1  g158(.A(G20), .B1(new_n294_), .B2(new_n186_), .ZN(new_n295_));
  AOI21_X1  g159(.A(new_n293_), .B1(new_n202_), .B2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g160(.A1(new_n285_), .A2(new_n289_), .A3(G190), .A4(new_n218_), .ZN(new_n297_));
  NAND4_X1  g161(.A1(new_n291_), .A2(new_n292_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  NAND2_X1  g162(.A1(new_n292_), .A2(new_n296_), .ZN(new_n299_));
  NAND2_X1  g163(.A1(new_n290_), .A2(new_n193_), .ZN(new_n300_));
  NAND4_X1  g164(.A1(new_n285_), .A2(new_n289_), .A3(new_n252_), .A4(new_n218_), .ZN(new_n301_));
  NAND3_X1  g165(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g166(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  OR4_X1    g167(.A1(new_n226_), .A2(new_n255_), .A3(new_n284_), .A4(new_n303_), .ZN(new_n304_));
  NAND3_X1  g168(.A1(new_n204_), .A2(new_n173_), .A3(G45), .ZN(new_n305_));
  OAI21_X1  g169(.A(KEYINPUT5), .B1(new_n179_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n307_));
  NOR3_X1   g171(.A1(new_n174_), .A2(G1), .A3(G41), .ZN(new_n308_));
  NAND4_X1  g172(.A1(new_n217_), .A2(new_n307_), .A3(new_n308_), .A4(G274), .ZN(new_n309_));
  NAND2_X1  g173(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g174(.A1(new_n184_), .A2(G257), .ZN(new_n311_));
  NAND3_X1  g175(.A1(new_n188_), .A2(G264), .A3(G1698), .ZN(new_n312_));
  NAND2_X1  g176(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g177(.A(G303), .ZN(new_n314_));
  NAND2_X1  g178(.A1(new_n314_), .A2(KEYINPUT16), .ZN(new_n315_));
  INV_X1    g179(.A(KEYINPUT16), .ZN(new_n316_));
  NAND2_X1  g180(.A1(new_n316_), .A2(G303), .ZN(new_n317_));
  AOI21_X1  g181(.A(new_n188_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g182(.A(new_n181_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g183(.A1(new_n181_), .A2(new_n308_), .ZN(new_n320_));
  NAND2_X1  g184(.A1(new_n320_), .A2(G270), .ZN(new_n321_));
  NAND4_X1  g185(.A1(new_n310_), .A2(G179), .A3(new_n319_), .A4(new_n321_), .ZN(new_n322_));
  INV_X1    g186(.A(KEYINPUT17), .ZN(new_n323_));
  NAND2_X1  g187(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g188(.A(KEYINPUT16), .B(G303), .ZN(new_n325_));
  OAI211_X1 g189(.A(new_n311_), .B(new_n312_), .C1(new_n325_), .C2(new_n188_), .ZN(new_n326_));
  AOI22_X1  g190(.A1(new_n326_), .A2(new_n181_), .B1(new_n320_), .B2(G270), .ZN(new_n327_));
  NAND4_X1  g191(.A1(new_n327_), .A2(KEYINPUT17), .A3(G179), .A4(new_n310_), .ZN(new_n328_));
  NAND2_X1  g192(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g193(.A1(new_n327_), .A2(new_n310_), .ZN(new_n330_));
  NAND2_X1  g194(.A1(new_n330_), .A2(G169), .ZN(new_n331_));
  NAND2_X1  g195(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g196(.A1(new_n204_), .A2(G33), .ZN(new_n333_));
  NAND4_X1  g197(.A1(new_n268_), .A2(G116), .A3(new_n269_), .A4(new_n333_), .ZN(new_n334_));
  NOR2_X1   g198(.A1(new_n198_), .A2(G116), .ZN(new_n335_));
  NOR2_X1   g199(.A1(new_n271_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g200(.A(G20), .B1(G33), .B2(G283), .ZN(new_n337_));
  OAI21_X1  g201(.A(new_n337_), .B1(G33), .B2(new_n286_), .ZN(new_n338_));
  AOI22_X1  g202(.A1(new_n336_), .A2(new_n338_), .B1(new_n276_), .B2(new_n335_), .ZN(new_n339_));
  NAND2_X1  g203(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g204(.A1(new_n332_), .A2(KEYINPUT18), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g205(.A(KEYINPUT18), .ZN(new_n342_));
  AOI22_X1  g206(.A1(new_n324_), .A2(new_n328_), .B1(G169), .B2(new_n330_), .ZN(new_n343_));
  INV_X1    g207(.A(new_n340_), .ZN(new_n344_));
  OAI21_X1  g208(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g209(.A(new_n340_), .B1(G200), .B2(new_n330_), .ZN(new_n346_));
  OAI21_X1  g210(.A(new_n346_), .B1(new_n236_), .B2(new_n330_), .ZN(new_n347_));
  NAND3_X1  g211(.A1(new_n341_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g212(.A(KEYINPUT8), .ZN(new_n349_));
  NAND3_X1  g213(.A1(new_n188_), .A2(G250), .A3(G1698), .ZN(new_n350_));
  NAND2_X1  g214(.A1(new_n350_), .A2(KEYINPUT3), .ZN(new_n351_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n352_));
  NAND4_X1  g216(.A1(new_n352_), .A2(new_n188_), .A3(G250), .A4(G1698), .ZN(new_n353_));
  NAND2_X1  g217(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  AOI22_X1  g218(.A1(new_n184_), .A2(G244), .B1(G33), .B2(G283), .ZN(new_n355_));
  NAND2_X1  g219(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g220(.A1(new_n356_), .A2(KEYINPUT4), .ZN(new_n357_));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n358_));
  NAND3_X1  g222(.A1(new_n354_), .A2(new_n358_), .A3(new_n355_), .ZN(new_n359_));
  AOI21_X1  g223(.A(new_n217_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n361_));
  NAND2_X1  g225(.A1(new_n217_), .A2(new_n305_), .ZN(new_n362_));
  INV_X1    g226(.A(G257), .ZN(new_n363_));
  OAI21_X1  g227(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g228(.A1(new_n217_), .A2(KEYINPUT6), .A3(G257), .A4(new_n305_), .ZN(new_n365_));
  NAND2_X1  g229(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g230(.A1(new_n366_), .A2(new_n310_), .ZN(new_n367_));
  OAI21_X1  g231(.A(new_n349_), .B1(new_n360_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g232(.A(new_n359_), .ZN(new_n369_));
  AOI21_X1  g233(.A(new_n358_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n370_));
  OAI21_X1  g234(.A(new_n181_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  AOI22_X1  g235(.A1(new_n364_), .A2(new_n365_), .B1(new_n309_), .B2(new_n306_), .ZN(new_n372_));
  NAND3_X1  g236(.A1(new_n371_), .A2(KEYINPUT8), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g237(.A(G20), .B1(G97), .B2(G107), .ZN(new_n374_));
  INV_X1    g238(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g239(.A(new_n375_), .B1(new_n286_), .B2(new_n168_), .ZN(new_n376_));
  INV_X1    g240(.A(G77), .ZN(new_n377_));
  OAI211_X1 g241(.A(new_n261_), .B(new_n198_), .C1(G33), .C2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g242(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n380_));
  NAND2_X1  g244(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g245(.A1(new_n376_), .A2(KEYINPUT7), .A3(new_n378_), .ZN(new_n382_));
  NAND3_X1  g246(.A1(new_n381_), .A2(new_n202_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g247(.A(new_n286_), .B1(new_n204_), .B2(G33), .ZN(new_n384_));
  AOI22_X1  g248(.A1(new_n209_), .A2(new_n384_), .B1(new_n286_), .B2(new_n206_), .ZN(new_n385_));
  AOI21_X1  g249(.A(new_n252_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g250(.A1(new_n368_), .A2(new_n373_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g251(.A1(new_n383_), .A2(new_n385_), .ZN(new_n388_));
  OAI211_X1 g252(.A(new_n388_), .B(G169), .C1(new_n360_), .C2(new_n367_), .ZN(new_n389_));
  AND2_X1   g253(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OR3_X1    g254(.A1(new_n174_), .A2(G1), .A3(G274), .ZN(new_n391_));
  INV_X1    g255(.A(G250), .ZN(new_n392_));
  OAI21_X1  g256(.A(new_n392_), .B1(new_n174_), .B2(G1), .ZN(new_n393_));
  NAND3_X1  g257(.A1(new_n391_), .A2(new_n217_), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g258(.A1(new_n188_), .A2(new_n230_), .A3(G238), .ZN(new_n395_));
  NAND3_X1  g259(.A1(new_n188_), .A2(G244), .A3(G1698), .ZN(new_n396_));
  NAND2_X1  g260(.A1(G33), .A2(G116), .ZN(new_n397_));
  NAND3_X1  g261(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  AND3_X1   g262(.A1(new_n398_), .A2(KEYINPUT14), .A3(new_n181_), .ZN(new_n399_));
  AOI21_X1  g263(.A(KEYINPUT14), .B1(new_n398_), .B2(new_n181_), .ZN(new_n400_));
  OAI211_X1 g264(.A(G190), .B(new_n394_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g265(.A(KEYINPUT13), .ZN(new_n402_));
  OAI21_X1  g266(.A(new_n402_), .B1(new_n199_), .B2(new_n286_), .ZN(new_n403_));
  NAND4_X1  g267(.A1(new_n198_), .A2(KEYINPUT13), .A3(G33), .A4(G97), .ZN(new_n404_));
  NAND2_X1  g268(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g269(.A(G87), .ZN(new_n406_));
  NAND3_X1  g270(.A1(new_n406_), .A2(new_n286_), .A3(new_n168_), .ZN(new_n407_));
  AOI22_X1  g271(.A1(new_n407_), .A2(G20), .B1(G68), .B2(new_n196_), .ZN(new_n408_));
  AOI21_X1  g272(.A(new_n271_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g273(.A1(new_n333_), .A2(G87), .ZN(new_n410_));
  OAI22_X1  g274(.A1(new_n208_), .A2(new_n410_), .B1(G87), .B2(new_n205_), .ZN(new_n411_));
  NOR2_X1   g275(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g276(.A1(new_n401_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g277(.A1(new_n398_), .A2(new_n181_), .ZN(new_n414_));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n415_));
  NAND2_X1  g279(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g280(.A1(new_n398_), .A2(KEYINPUT14), .A3(new_n181_), .ZN(new_n417_));
  NAND2_X1  g281(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g282(.A(new_n223_), .B1(new_n418_), .B2(new_n394_), .ZN(new_n419_));
  NOR2_X1   g283(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g284(.A(KEYINPUT15), .ZN(new_n421_));
  INV_X1    g285(.A(new_n394_), .ZN(new_n422_));
  AOI21_X1  g286(.A(new_n422_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n423_));
  OAI21_X1  g287(.A(new_n421_), .B1(new_n423_), .B2(new_n193_), .ZN(new_n424_));
  NAND2_X1  g288(.A1(new_n423_), .A2(G179), .ZN(new_n425_));
  OAI21_X1  g289(.A(new_n394_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n426_));
  NAND3_X1  g290(.A1(new_n426_), .A2(KEYINPUT15), .A3(G169), .ZN(new_n427_));
  NAND3_X1  g291(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g292(.A(new_n412_), .ZN(new_n429_));
  AOI21_X1  g293(.A(new_n420_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g294(.A(G200), .B1(new_n360_), .B2(new_n367_), .ZN(new_n431_));
  INV_X1    g295(.A(new_n388_), .ZN(new_n432_));
  NAND3_X1  g296(.A1(new_n371_), .A2(G190), .A3(new_n372_), .ZN(new_n433_));
  NAND3_X1  g297(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g298(.A1(new_n168_), .A2(G20), .ZN(new_n435_));
  XNOR2_X1  g299(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  NAND2_X1  g300(.A1(new_n188_), .A2(G87), .ZN(new_n437_));
  AOI21_X1  g301(.A(G20), .B1(new_n437_), .B2(new_n397_), .ZN(new_n438_));
  OAI21_X1  g302(.A(new_n202_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g303(.A1(new_n209_), .A2(G107), .A3(new_n333_), .ZN(new_n440_));
  NAND2_X1  g304(.A1(new_n206_), .A2(new_n168_), .ZN(new_n441_));
  NAND3_X1  g305(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g306(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g307(.A1(G33), .A2(G294), .ZN(new_n444_));
  OAI221_X1 g308(.A(new_n444_), .B1(new_n189_), .B2(new_n363_), .C1(new_n392_), .C2(new_n231_), .ZN(new_n445_));
  AOI22_X1  g309(.A1(new_n445_), .A2(new_n181_), .B1(new_n320_), .B2(G264), .ZN(new_n446_));
  NAND2_X1  g310(.A1(new_n446_), .A2(new_n310_), .ZN(new_n447_));
  AOI21_X1  g311(.A(new_n443_), .B1(new_n193_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g312(.A1(new_n446_), .A2(new_n310_), .ZN(new_n449_));
  NAND2_X1  g313(.A1(new_n449_), .A2(new_n252_), .ZN(new_n450_));
  AOI21_X1  g314(.A(new_n442_), .B1(new_n449_), .B2(G190), .ZN(new_n451_));
  NAND2_X1  g315(.A1(new_n447_), .A2(G200), .ZN(new_n452_));
  AOI22_X1  g316(.A1(new_n448_), .A2(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g317(.A1(new_n390_), .A2(new_n430_), .A3(new_n434_), .A4(new_n453_), .ZN(new_n454_));
  NOR3_X1   g318(.A1(new_n304_), .A2(new_n348_), .A3(new_n454_), .ZN(G372));
  INV_X1    g319(.A(new_n302_), .ZN(new_n456_));
  NAND2_X1  g320(.A1(new_n254_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g321(.A1(new_n457_), .A2(new_n226_), .ZN(new_n458_));
  XNOR2_X1  g322(.A(new_n458_), .B(KEYINPUT20), .ZN(new_n459_));
  AOI211_X1 g323(.A(new_n303_), .B(new_n283_), .C1(new_n240_), .C2(new_n249_), .ZN(new_n460_));
  NAND2_X1  g324(.A1(new_n251_), .A2(new_n253_), .ZN(new_n461_));
  INV_X1    g325(.A(new_n461_), .ZN(new_n462_));
  OAI211_X1 g326(.A(new_n225_), .B(new_n220_), .C1(new_n460_), .C2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g327(.A1(new_n459_), .A2(new_n213_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g328(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g329(.A(new_n193_), .B1(new_n418_), .B2(new_n394_), .ZN(new_n466_));
  AOI22_X1  g330(.A1(new_n466_), .A2(KEYINPUT15), .B1(G179), .B2(new_n423_), .ZN(new_n467_));
  AOI21_X1  g331(.A(new_n412_), .B1(new_n467_), .B2(new_n424_), .ZN(new_n468_));
  NAND2_X1  g332(.A1(new_n387_), .A2(new_n389_), .ZN(new_n469_));
  INV_X1    g333(.A(new_n420_), .ZN(new_n470_));
  AOI21_X1  g334(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g335(.A1(new_n430_), .A2(new_n387_), .A3(new_n389_), .A4(new_n434_), .ZN(new_n472_));
  NAND2_X1  g336(.A1(new_n447_), .A2(new_n193_), .ZN(new_n473_));
  AND3_X1   g337(.A1(new_n450_), .A2(new_n442_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g338(.A(new_n344_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n475_));
  OAI211_X1 g339(.A(new_n452_), .B(new_n443_), .C1(new_n236_), .C2(new_n447_), .ZN(new_n476_));
  AOI21_X1  g340(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g341(.A(new_n471_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g342(.A(new_n478_), .ZN(new_n479_));
  OAI21_X1  g343(.A(new_n465_), .B1(new_n304_), .B2(new_n479_), .ZN(G369));
  NAND3_X1  g344(.A1(new_n276_), .A2(new_n198_), .A3(G213), .ZN(new_n481_));
  INV_X1    g345(.A(G343), .ZN(new_n482_));
  NOR2_X1   g346(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g347(.A1(new_n442_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g348(.A1(new_n453_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g349(.A1(new_n474_), .A2(new_n442_), .A3(new_n483_), .ZN(new_n486_));
  NAND2_X1  g350(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND3_X1   g351(.A1(new_n341_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n488_));
  INV_X1    g352(.A(new_n483_), .ZN(new_n489_));
  NOR2_X1   g353(.A1(new_n344_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g354(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g355(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n493_));
  NAND2_X1  g357(.A1(new_n341_), .A2(new_n345_), .ZN(new_n494_));
  NAND2_X1  g358(.A1(new_n494_), .A2(new_n490_), .ZN(new_n495_));
  AND3_X1   g359(.A1(new_n492_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g360(.A(new_n493_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n497_));
  OAI211_X1 g361(.A(G330), .B(new_n487_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g362(.A(new_n483_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n499_));
  AOI22_X1  g363(.A1(new_n487_), .A2(new_n499_), .B1(new_n474_), .B2(new_n489_), .ZN(new_n500_));
  NAND2_X1  g364(.A1(new_n498_), .A2(new_n500_), .ZN(G399));
  NOR2_X1   g365(.A1(new_n144_), .A2(G41), .ZN(new_n502_));
  INV_X1    g366(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g367(.A1(new_n407_), .A2(G116), .ZN(new_n504_));
  NAND3_X1  g368(.A1(new_n503_), .A2(G1), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g369(.A(G330), .ZN(new_n506_));
  NAND3_X1  g370(.A1(new_n434_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n507_));
  NAND2_X1  g371(.A1(new_n427_), .A2(new_n425_), .ZN(new_n508_));
  AOI21_X1  g372(.A(KEYINPUT15), .B1(new_n426_), .B2(G169), .ZN(new_n509_));
  OAI21_X1  g373(.A(new_n429_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g374(.A1(new_n510_), .A2(new_n470_), .ZN(new_n511_));
  NOR2_X1   g375(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND4_X1  g376(.A1(new_n488_), .A2(new_n512_), .A3(new_n453_), .A4(new_n489_), .ZN(new_n513_));
  NAND2_X1  g377(.A1(new_n368_), .A2(new_n373_), .ZN(new_n514_));
  NOR2_X1   g378(.A1(new_n449_), .A2(G179), .ZN(new_n515_));
  NAND4_X1  g379(.A1(new_n514_), .A2(new_n330_), .A3(new_n426_), .A4(new_n515_), .ZN(new_n516_));
  INV_X1    g380(.A(new_n329_), .ZN(new_n517_));
  NOR2_X1   g381(.A1(new_n360_), .A2(new_n367_), .ZN(new_n518_));
  NAND4_X1  g382(.A1(new_n517_), .A2(new_n423_), .A3(new_n518_), .A4(new_n449_), .ZN(new_n519_));
  AOI21_X1  g383(.A(new_n489_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g384(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g385(.A(new_n506_), .B1(new_n513_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g386(.A1(new_n332_), .A2(new_n476_), .A3(new_n340_), .ZN(new_n523_));
  INV_X1    g387(.A(new_n474_), .ZN(new_n524_));
  NAND2_X1  g388(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AND3_X1   g389(.A1(new_n434_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n526_));
  NAND3_X1  g390(.A1(new_n525_), .A2(new_n526_), .A3(new_n430_), .ZN(new_n527_));
  AOI21_X1  g391(.A(new_n483_), .B1(new_n527_), .B2(new_n471_), .ZN(new_n528_));
  NOR2_X1   g392(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  OAI221_X1 g393(.A(new_n505_), .B1(new_n146_), .B2(new_n503_), .C1(new_n529_), .C2(G1), .ZN(G364));
  NOR2_X1   g394(.A1(new_n275_), .A2(G20), .ZN(new_n531_));
  AOI21_X1  g395(.A(new_n204_), .B1(new_n531_), .B2(G45), .ZN(new_n532_));
  INV_X1    g396(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g397(.A1(new_n502_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g398(.A1(new_n143_), .A2(new_n188_), .ZN(new_n535_));
  INV_X1    g399(.A(G355), .ZN(new_n536_));
  OAI22_X1  g400(.A1(new_n535_), .A2(new_n536_), .B1(G116), .B2(new_n143_), .ZN(new_n537_));
  NAND2_X1  g401(.A1(new_n165_), .A2(G45), .ZN(new_n538_));
  NAND2_X1  g402(.A1(new_n143_), .A2(G33), .ZN(new_n539_));
  INV_X1    g403(.A(new_n146_), .ZN(new_n540_));
  AOI21_X1  g404(.A(new_n539_), .B1(new_n540_), .B2(new_n174_), .ZN(new_n541_));
  AOI21_X1  g405(.A(new_n537_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g406(.A1(G13), .A2(G33), .ZN(new_n543_));
  XOR2_X1   g407(.A(new_n543_), .B(KEYINPUT28), .Z(new_n544_));
  NOR2_X1   g408(.A1(new_n544_), .A2(G20), .ZN(new_n545_));
  AOI21_X1  g409(.A(new_n178_), .B1(G20), .B2(new_n193_), .ZN(new_n546_));
  NOR2_X1   g410(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g411(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g412(.A(new_n534_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g413(.A1(new_n236_), .A2(G20), .ZN(new_n550_));
  OR2_X1    g414(.A1(new_n550_), .A2(KEYINPUT22), .ZN(new_n551_));
  NAND2_X1  g415(.A1(new_n550_), .A2(KEYINPUT22), .ZN(new_n552_));
  NAND2_X1  g416(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g417(.A1(new_n198_), .A2(new_n252_), .A3(G200), .ZN(new_n554_));
  NAND2_X1  g418(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR3_X1   g419(.A1(new_n198_), .A2(new_n252_), .A3(new_n223_), .ZN(new_n556_));
  NAND2_X1  g420(.A1(new_n556_), .A2(G190), .ZN(new_n557_));
  OAI22_X1  g421(.A1(new_n555_), .A2(new_n137_), .B1(new_n203_), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g422(.A(new_n558_), .B(KEYINPUT23), .ZN(new_n559_));
  NAND2_X1  g423(.A1(new_n554_), .A2(new_n236_), .ZN(new_n560_));
  OAI21_X1  g424(.A(G20), .B1(G179), .B2(G200), .ZN(new_n561_));
  NAND2_X1  g425(.A1(new_n550_), .A2(new_n561_), .ZN(new_n562_));
  OAI22_X1  g426(.A1(new_n560_), .A2(new_n377_), .B1(new_n286_), .B2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g427(.A1(new_n198_), .A2(G179), .ZN(new_n564_));
  NAND3_X1  g428(.A1(new_n564_), .A2(G190), .A3(G200), .ZN(new_n565_));
  NOR2_X1   g429(.A1(new_n565_), .A2(new_n406_), .ZN(new_n566_));
  NOR2_X1   g430(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g431(.A1(new_n564_), .A2(new_n236_), .A3(G200), .ZN(new_n568_));
  NAND3_X1  g432(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n569_));
  OAI221_X1 g433(.A(new_n188_), .B1(new_n168_), .B2(new_n568_), .C1(new_n569_), .C2(new_n138_), .ZN(new_n570_));
  NAND3_X1  g434(.A1(new_n551_), .A2(new_n552_), .A3(new_n561_), .ZN(new_n571_));
  INV_X1    g435(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g436(.A(new_n570_), .B1(G159), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g437(.A1(new_n559_), .A2(new_n567_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g438(.A(G283), .ZN(new_n575_));
  NOR2_X1   g439(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g440(.A(new_n576_), .B(KEYINPUT25), .ZN(new_n577_));
  INV_X1    g441(.A(G322), .ZN(new_n578_));
  INV_X1    g442(.A(G317), .ZN(new_n579_));
  OAI22_X1  g443(.A1(new_n555_), .A2(new_n578_), .B1(new_n579_), .B2(new_n569_), .ZN(new_n580_));
  INV_X1    g444(.A(G326), .ZN(new_n581_));
  INV_X1    g445(.A(G294), .ZN(new_n582_));
  OAI22_X1  g446(.A1(new_n557_), .A2(new_n581_), .B1(new_n582_), .B2(new_n562_), .ZN(new_n583_));
  INV_X1    g447(.A(G311), .ZN(new_n584_));
  OAI22_X1  g448(.A1(new_n560_), .A2(new_n584_), .B1(new_n565_), .B2(new_n325_), .ZN(new_n585_));
  NOR3_X1   g449(.A1(new_n580_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g450(.A(new_n586_), .B(KEYINPUT24), .ZN(new_n587_));
  AOI211_X1 g451(.A(new_n577_), .B(new_n587_), .C1(G329), .C2(new_n572_), .ZN(new_n588_));
  INV_X1    g452(.A(KEYINPUT26), .ZN(new_n589_));
  AND2_X1   g453(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g454(.A(G33), .B1(new_n588_), .B2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g455(.A(new_n574_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g456(.A1(new_n592_), .A2(KEYINPUT27), .ZN(new_n593_));
  INV_X1    g457(.A(new_n546_), .ZN(new_n594_));
  AOI21_X1  g458(.A(new_n594_), .B1(new_n592_), .B2(KEYINPUT27), .ZN(new_n595_));
  AOI21_X1  g459(.A(new_n549_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g460(.A1(new_n496_), .A2(new_n497_), .ZN(new_n597_));
  NAND2_X1  g461(.A1(new_n597_), .A2(new_n545_), .ZN(new_n598_));
  NAND2_X1  g462(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g463(.A1(new_n492_), .A2(new_n495_), .ZN(new_n600_));
  NAND2_X1  g464(.A1(new_n600_), .A2(KEYINPUT21), .ZN(new_n601_));
  NAND3_X1  g465(.A1(new_n492_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n602_));
  AOI21_X1  g466(.A(new_n506_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g467(.A1(new_n603_), .A2(new_n534_), .ZN(new_n604_));
  NAND2_X1  g468(.A1(new_n597_), .A2(new_n506_), .ZN(new_n605_));
  NAND2_X1  g469(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g470(.A1(new_n599_), .A2(new_n606_), .ZN(G396));
  XNOR2_X1  g471(.A(new_n522_), .B(KEYINPUT29), .ZN(new_n608_));
  NAND2_X1  g472(.A1(new_n478_), .A2(new_n489_), .ZN(new_n609_));
  NAND2_X1  g473(.A1(new_n281_), .A2(new_n483_), .ZN(new_n610_));
  NAND3_X1  g474(.A1(new_n279_), .A2(new_n283_), .A3(new_n610_), .ZN(new_n611_));
  NAND4_X1  g475(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .A4(new_n483_), .ZN(new_n612_));
  NAND2_X1  g476(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g477(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g478(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g479(.A1(new_n478_), .A2(new_n489_), .A3(new_n613_), .ZN(new_n616_));
  NAND2_X1  g480(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g481(.A(new_n534_), .B1(new_n608_), .B2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g482(.A(new_n618_), .B1(new_n617_), .B2(new_n608_), .ZN(new_n619_));
  OR2_X1    g483(.A1(new_n546_), .A2(new_n543_), .ZN(new_n620_));
  OAI21_X1  g484(.A(new_n534_), .B1(new_n620_), .B2(G77), .ZN(new_n621_));
  NOR2_X1   g485(.A1(new_n568_), .A2(new_n406_), .ZN(new_n622_));
  INV_X1    g486(.A(new_n560_), .ZN(new_n623_));
  AOI21_X1  g487(.A(new_n622_), .B1(G116), .B2(new_n623_), .ZN(new_n624_));
  OAI221_X1 g488(.A(new_n624_), .B1(new_n168_), .B2(new_n565_), .C1(new_n314_), .C2(new_n557_), .ZN(new_n625_));
  INV_X1    g489(.A(new_n569_), .ZN(new_n626_));
  AOI22_X1  g490(.A1(G311), .A2(new_n572_), .B1(new_n626_), .B2(G283), .ZN(new_n627_));
  INV_X1    g491(.A(new_n562_), .ZN(new_n628_));
  AOI21_X1  g492(.A(new_n188_), .B1(new_n628_), .B2(G97), .ZN(new_n629_));
  OAI211_X1 g493(.A(new_n627_), .B(new_n629_), .C1(new_n582_), .C2(new_n555_), .ZN(new_n630_));
  OAI21_X1  g494(.A(new_n188_), .B1(new_n565_), .B2(new_n203_), .ZN(new_n631_));
  AOI21_X1  g495(.A(new_n631_), .B1(new_n572_), .B2(G132), .ZN(new_n632_));
  INV_X1    g496(.A(G143), .ZN(new_n633_));
  INV_X1    g497(.A(G150), .ZN(new_n634_));
  OAI221_X1 g498(.A(new_n632_), .B1(new_n633_), .B2(new_n555_), .C1(new_n634_), .C2(new_n569_), .ZN(new_n635_));
  AOI22_X1  g499(.A1(new_n623_), .A2(G159), .B1(G58), .B2(new_n628_), .ZN(new_n636_));
  INV_X1    g500(.A(G137), .ZN(new_n637_));
  OAI221_X1 g501(.A(new_n636_), .B1(new_n138_), .B2(new_n568_), .C1(new_n637_), .C2(new_n557_), .ZN(new_n638_));
  OAI22_X1  g502(.A1(new_n625_), .A2(new_n630_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  OR2_X1    g503(.A1(new_n639_), .A2(KEYINPUT30), .ZN(new_n640_));
  AOI21_X1  g504(.A(new_n594_), .B1(new_n639_), .B2(KEYINPUT30), .ZN(new_n641_));
  AOI21_X1  g505(.A(new_n621_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g506(.A(new_n642_), .B1(new_n544_), .B2(new_n613_), .ZN(new_n643_));
  AND2_X1   g507(.A1(new_n619_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g508(.A(new_n644_), .ZN(G384));
  NOR2_X1   g509(.A1(new_n531_), .A2(new_n204_), .ZN(new_n646_));
  NOR2_X1   g510(.A1(new_n609_), .A2(new_n304_), .ZN(new_n647_));
  OR2_X1    g511(.A1(new_n464_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g512(.A(new_n481_), .ZN(new_n649_));
  NAND2_X1  g513(.A1(new_n248_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g514(.A(new_n650_), .ZN(new_n651_));
  AND3_X1   g515(.A1(new_n251_), .A2(new_n253_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g516(.A(new_n652_), .B1(new_n254_), .B2(new_n650_), .ZN(new_n653_));
  NAND2_X1  g517(.A1(new_n456_), .A2(new_n489_), .ZN(new_n654_));
  OAI22_X1  g518(.A1(new_n653_), .A2(new_n654_), .B1(new_n461_), .B2(new_n649_), .ZN(new_n655_));
  INV_X1    g519(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g520(.A1(new_n254_), .A2(new_n650_), .ZN(new_n657_));
  INV_X1    g521(.A(new_n652_), .ZN(new_n658_));
  NAND2_X1  g522(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g523(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .A4(new_n483_), .ZN(new_n660_));
  XNOR2_X1  g524(.A(new_n660_), .B(KEYINPUT31), .ZN(new_n661_));
  INV_X1    g525(.A(KEYINPUT32), .ZN(new_n662_));
  NAND2_X1  g526(.A1(new_n299_), .A2(new_n483_), .ZN(new_n663_));
  NAND4_X1  g527(.A1(new_n298_), .A2(new_n302_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n664_));
  NAND3_X1  g528(.A1(new_n298_), .A2(new_n302_), .A3(new_n663_), .ZN(new_n665_));
  NAND2_X1  g529(.A1(new_n665_), .A2(KEYINPUT32), .ZN(new_n666_));
  NAND3_X1  g530(.A1(new_n661_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  NOR2_X1   g531(.A1(new_n283_), .A2(new_n483_), .ZN(new_n668_));
  NAND3_X1  g532(.A1(new_n659_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g533(.A1(new_n656_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g534(.A(new_n667_), .ZN(new_n671_));
  NAND4_X1  g535(.A1(new_n478_), .A2(new_n489_), .A3(new_n613_), .A4(new_n659_), .ZN(new_n672_));
  AOI21_X1  g536(.A(new_n671_), .B1(new_n672_), .B2(KEYINPUT33), .ZN(new_n673_));
  INV_X1    g537(.A(KEYINPUT33), .ZN(new_n674_));
  NAND4_X1  g538(.A1(new_n528_), .A2(new_n674_), .A3(new_n613_), .A4(new_n659_), .ZN(new_n675_));
  AOI21_X1  g539(.A(new_n670_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g540(.A(new_n648_), .B(new_n676_), .ZN(new_n677_));
  NAND3_X1  g541(.A1(new_n659_), .A2(new_n667_), .A3(new_n613_), .ZN(new_n678_));
  AND2_X1   g542(.A1(new_n304_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g543(.A(new_n522_), .ZN(new_n680_));
  INV_X1    g544(.A(new_n678_), .ZN(new_n681_));
  AOI21_X1  g545(.A(new_n304_), .B1(new_n521_), .B2(new_n513_), .ZN(new_n682_));
  AOI211_X1 g546(.A(new_n679_), .B(new_n680_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g547(.A(new_n646_), .B1(new_n677_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g548(.A(new_n684_), .B1(new_n677_), .B2(new_n683_), .ZN(new_n685_));
  INV_X1    g549(.A(G116), .ZN(new_n686_));
  NOR3_X1   g550(.A1(new_n376_), .A2(new_n686_), .A3(new_n178_), .ZN(new_n687_));
  NAND2_X1  g551(.A1(new_n244_), .A2(G77), .ZN(new_n688_));
  OAI22_X1  g552(.A1(new_n146_), .A2(new_n688_), .B1(G50), .B2(new_n138_), .ZN(new_n689_));
  NOR2_X1   g553(.A1(new_n204_), .A2(G13), .ZN(new_n690_));
  AOI21_X1  g554(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g555(.A1(new_n685_), .A2(new_n691_), .ZN(G367));
  INV_X1    g556(.A(new_n529_), .ZN(new_n693_));
  NAND2_X1  g557(.A1(new_n388_), .A2(new_n483_), .ZN(new_n694_));
  NAND2_X1  g558(.A1(new_n526_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g559(.A1(new_n469_), .A2(new_n388_), .A3(new_n483_), .ZN(new_n696_));
  AND2_X1   g560(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g561(.A(KEYINPUT35), .ZN(new_n698_));
  NAND2_X1  g562(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g563(.A(new_n500_), .ZN(new_n700_));
  NAND2_X1  g564(.A1(new_n695_), .A2(new_n696_), .ZN(new_n701_));
  NAND2_X1  g565(.A1(new_n701_), .A2(KEYINPUT35), .ZN(new_n702_));
  NAND3_X1  g566(.A1(new_n699_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  NAND3_X1  g567(.A1(new_n500_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n704_));
  NAND2_X1  g568(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g569(.A1(new_n705_), .A2(new_n487_), .A3(new_n603_), .ZN(new_n706_));
  NAND3_X1  g570(.A1(new_n498_), .A2(new_n704_), .A3(new_n703_), .ZN(new_n707_));
  NAND2_X1  g571(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g572(.A(new_n487_), .B(new_n499_), .Z(new_n709_));
  INV_X1    g573(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g574(.A(new_n710_), .B1(new_n597_), .B2(new_n506_), .ZN(new_n711_));
  NAND2_X1  g575(.A1(new_n603_), .A2(new_n709_), .ZN(new_n712_));
  AND2_X1   g576(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g577(.A(new_n693_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g578(.A(new_n532_), .B1(new_n714_), .B2(new_n503_), .ZN(new_n715_));
  OAI22_X1  g579(.A1(new_n500_), .A2(new_n697_), .B1(new_n390_), .B2(new_n483_), .ZN(new_n716_));
  NAND2_X1  g580(.A1(new_n716_), .A2(KEYINPUT34), .ZN(new_n717_));
  OAI21_X1  g581(.A(new_n430_), .B1(new_n412_), .B2(new_n489_), .ZN(new_n718_));
  OAI21_X1  g582(.A(new_n718_), .B1(new_n510_), .B2(new_n489_), .ZN(new_n719_));
  NAND2_X1  g583(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND4_X1  g584(.A1(new_n720_), .A2(new_n487_), .A3(new_n603_), .A4(new_n701_), .ZN(new_n721_));
  OAI211_X1 g585(.A(new_n719_), .B(new_n717_), .C1(new_n498_), .C2(new_n697_), .ZN(new_n722_));
  NOR2_X1   g586(.A1(new_n716_), .A2(KEYINPUT34), .ZN(new_n723_));
  AND3_X1   g587(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g588(.A(new_n723_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n725_));
  NOR2_X1   g589(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g590(.A1(new_n715_), .A2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g591(.A1(new_n158_), .A2(new_n539_), .ZN(new_n728_));
  OAI21_X1  g592(.A(new_n547_), .B1(new_n406_), .B2(new_n143_), .ZN(new_n729_));
  OAI21_X1  g593(.A(new_n534_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g594(.A(new_n188_), .B1(new_n565_), .B2(new_n137_), .ZN(new_n731_));
  AOI21_X1  g595(.A(new_n731_), .B1(new_n572_), .B2(G137), .ZN(new_n732_));
  INV_X1    g596(.A(G159), .ZN(new_n733_));
  OAI221_X1 g597(.A(new_n732_), .B1(new_n634_), .B2(new_n555_), .C1(new_n733_), .C2(new_n569_), .ZN(new_n734_));
  OAI22_X1  g598(.A1(new_n557_), .A2(new_n633_), .B1(new_n138_), .B2(new_n562_), .ZN(new_n735_));
  OAI22_X1  g599(.A1(new_n560_), .A2(new_n203_), .B1(new_n568_), .B2(new_n377_), .ZN(new_n736_));
  NOR3_X1   g600(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  OR2_X1    g601(.A1(new_n737_), .A2(KEYINPUT36), .ZN(new_n738_));
  NAND2_X1  g602(.A1(new_n737_), .A2(KEYINPUT36), .ZN(new_n739_));
  OAI22_X1  g603(.A1(new_n557_), .A2(new_n584_), .B1(new_n168_), .B2(new_n562_), .ZN(new_n740_));
  OAI221_X1 g604(.A(G33), .B1(new_n286_), .B2(new_n568_), .C1(new_n555_), .C2(new_n314_), .ZN(new_n741_));
  OAI22_X1  g605(.A1(new_n560_), .A2(new_n575_), .B1(new_n565_), .B2(new_n686_), .ZN(new_n742_));
  XNOR2_X1  g606(.A(KEYINPUT37), .B(G294), .ZN(new_n743_));
  OAI22_X1  g607(.A1(new_n569_), .A2(new_n743_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n744_));
  OR4_X1    g608(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .A4(new_n744_), .ZN(new_n745_));
  NAND3_X1  g609(.A1(new_n738_), .A2(new_n739_), .A3(new_n745_), .ZN(new_n746_));
  AOI21_X1  g610(.A(new_n730_), .B1(new_n746_), .B2(new_n546_), .ZN(new_n747_));
  INV_X1    g611(.A(new_n545_), .ZN(new_n748_));
  OAI21_X1  g612(.A(new_n747_), .B1(new_n719_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g613(.A1(new_n727_), .A2(new_n749_), .ZN(G387));
  NAND2_X1  g614(.A1(new_n711_), .A2(new_n712_), .ZN(new_n751_));
  NAND2_X1  g615(.A1(new_n751_), .A2(new_n693_), .ZN(new_n752_));
  NAND3_X1  g616(.A1(new_n711_), .A2(new_n712_), .A3(new_n529_), .ZN(new_n753_));
  NAND3_X1  g617(.A1(new_n752_), .A2(new_n502_), .A3(new_n753_), .ZN(new_n754_));
  NAND3_X1  g618(.A1(new_n485_), .A2(new_n486_), .A3(new_n545_), .ZN(new_n755_));
  OAI21_X1  g619(.A(new_n174_), .B1(new_n138_), .B2(new_n377_), .ZN(new_n756_));
  NOR3_X1   g620(.A1(new_n756_), .A2(G50), .A3(new_n137_), .ZN(new_n757_));
  AOI21_X1  g621(.A(new_n539_), .B1(new_n757_), .B2(new_n504_), .ZN(new_n758_));
  OAI21_X1  g622(.A(new_n758_), .B1(new_n161_), .B2(new_n174_), .ZN(new_n759_));
  XNOR2_X1  g623(.A(new_n759_), .B(KEYINPUT40), .ZN(new_n760_));
  OAI22_X1  g624(.A1(new_n504_), .A2(new_n535_), .B1(G107), .B2(new_n143_), .ZN(new_n761_));
  OAI21_X1  g625(.A(new_n547_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g626(.A1(new_n762_), .A2(new_n534_), .ZN(new_n763_));
  OAI221_X1 g627(.A(G33), .B1(new_n575_), .B2(new_n562_), .C1(new_n569_), .C2(new_n584_), .ZN(new_n764_));
  INV_X1    g628(.A(new_n555_), .ZN(new_n765_));
  AOI21_X1  g629(.A(new_n764_), .B1(G317), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g630(.A1(new_n571_), .A2(new_n581_), .ZN(new_n767_));
  XNOR2_X1  g631(.A(new_n767_), .B(KEYINPUT39), .ZN(new_n768_));
  OAI22_X1  g632(.A1(new_n557_), .A2(new_n578_), .B1(new_n565_), .B2(new_n743_), .ZN(new_n769_));
  OAI22_X1  g633(.A1(new_n560_), .A2(new_n325_), .B1(new_n568_), .B2(new_n686_), .ZN(new_n770_));
  NOR2_X1   g634(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g635(.A1(new_n766_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  OAI221_X1 g636(.A(new_n188_), .B1(new_n286_), .B2(new_n568_), .C1(new_n569_), .C2(new_n137_), .ZN(new_n773_));
  AOI21_X1  g637(.A(new_n773_), .B1(G150), .B2(new_n572_), .ZN(new_n774_));
  NOR2_X1   g638(.A1(new_n562_), .A2(new_n406_), .ZN(new_n775_));
  NOR2_X1   g639(.A1(new_n565_), .A2(new_n377_), .ZN(new_n776_));
  AOI211_X1 g640(.A(new_n775_), .B(new_n776_), .C1(G68), .C2(new_n623_), .ZN(new_n777_));
  NAND2_X1  g641(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  OAI22_X1  g642(.A1(new_n555_), .A2(new_n203_), .B1(new_n733_), .B2(new_n557_), .ZN(new_n779_));
  XNOR2_X1  g643(.A(new_n779_), .B(KEYINPUT38), .ZN(new_n780_));
  OAI21_X1  g644(.A(new_n772_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g645(.A(new_n763_), .B1(new_n546_), .B2(new_n781_), .ZN(new_n782_));
  AOI22_X1  g646(.A1(new_n713_), .A2(new_n533_), .B1(new_n755_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g647(.A1(new_n754_), .A2(new_n783_), .ZN(G393));
  NAND2_X1  g648(.A1(new_n706_), .A2(KEYINPUT41), .ZN(new_n785_));
  NAND2_X1  g649(.A1(new_n785_), .A2(new_n753_), .ZN(new_n786_));
  AOI21_X1  g650(.A(new_n503_), .B1(new_n786_), .B2(new_n708_), .ZN(new_n787_));
  AND2_X1   g651(.A1(new_n706_), .A2(new_n707_), .ZN(new_n788_));
  NAND3_X1  g652(.A1(new_n788_), .A2(new_n753_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g653(.A1(new_n697_), .A2(new_n545_), .ZN(new_n790_));
  AND3_X1   g654(.A1(new_n171_), .A2(G33), .A3(new_n143_), .ZN(new_n791_));
  OAI21_X1  g655(.A(new_n547_), .B1(new_n286_), .B2(new_n143_), .ZN(new_n792_));
  OAI21_X1  g656(.A(new_n534_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  AOI211_X1 g657(.A(G33), .B(new_n622_), .C1(new_n765_), .C2(G159), .ZN(new_n794_));
  INV_X1    g658(.A(new_n557_), .ZN(new_n795_));
  AOI22_X1  g659(.A1(new_n795_), .A2(G150), .B1(new_n628_), .B2(G77), .ZN(new_n796_));
  INV_X1    g660(.A(new_n565_), .ZN(new_n797_));
  AOI22_X1  g661(.A1(new_n623_), .A2(G58), .B1(new_n797_), .B2(G68), .ZN(new_n798_));
  AOI22_X1  g662(.A1(G143), .A2(new_n572_), .B1(new_n626_), .B2(G50), .ZN(new_n799_));
  NAND4_X1  g663(.A1(new_n794_), .A2(new_n796_), .A3(new_n798_), .A4(new_n799_), .ZN(new_n800_));
  OAI22_X1  g664(.A1(new_n555_), .A2(new_n584_), .B1(new_n325_), .B2(new_n569_), .ZN(new_n801_));
  OAI22_X1  g665(.A1(new_n557_), .A2(new_n579_), .B1(new_n686_), .B2(new_n562_), .ZN(new_n802_));
  OAI22_X1  g666(.A1(new_n560_), .A2(new_n743_), .B1(new_n565_), .B2(new_n575_), .ZN(new_n803_));
  NOR3_X1   g667(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g668(.A(new_n804_), .B(KEYINPUT42), .ZN(new_n805_));
  OAI221_X1 g669(.A(G33), .B1(new_n168_), .B2(new_n568_), .C1(new_n571_), .C2(new_n578_), .ZN(new_n806_));
  OAI21_X1  g670(.A(new_n800_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g671(.A(new_n793_), .B1(new_n807_), .B2(new_n546_), .ZN(new_n808_));
  NAND2_X1  g672(.A1(new_n790_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g673(.A(KEYINPUT43), .B(new_n809_), .C1(new_n788_), .C2(new_n532_), .ZN(new_n810_));
  INV_X1    g674(.A(KEYINPUT43), .ZN(new_n811_));
  AOI21_X1  g675(.A(new_n532_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n812_));
  INV_X1    g676(.A(new_n809_), .ZN(new_n813_));
  OAI21_X1  g677(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI22_X1  g678(.A1(new_n787_), .A2(new_n789_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g679(.A(new_n815_), .ZN(G390));
  INV_X1    g680(.A(new_n668_), .ZN(new_n817_));
  NAND3_X1  g681(.A1(new_n616_), .A2(new_n667_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g682(.A1(new_n818_), .A2(new_n522_), .A3(new_n613_), .ZN(new_n819_));
  INV_X1    g683(.A(KEYINPUT46), .ZN(new_n820_));
  AOI211_X1 g684(.A(new_n820_), .B(new_n667_), .C1(new_n616_), .C2(new_n817_), .ZN(new_n821_));
  NOR2_X1   g685(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g686(.A(new_n668_), .B1(new_n528_), .B2(new_n613_), .ZN(new_n823_));
  OAI21_X1  g687(.A(new_n820_), .B1(new_n823_), .B2(new_n667_), .ZN(new_n824_));
  NAND2_X1  g688(.A1(new_n616_), .A2(new_n817_), .ZN(new_n825_));
  NAND2_X1  g689(.A1(new_n825_), .A2(new_n671_), .ZN(new_n826_));
  INV_X1    g690(.A(KEYINPUT47), .ZN(new_n827_));
  NAND3_X1  g691(.A1(new_n826_), .A2(new_n827_), .A3(new_n818_), .ZN(new_n828_));
  AOI21_X1  g692(.A(new_n667_), .B1(new_n616_), .B2(new_n817_), .ZN(new_n829_));
  AOI22_X1  g693(.A1(new_n829_), .A2(KEYINPUT47), .B1(new_n522_), .B2(new_n613_), .ZN(new_n830_));
  AOI22_X1  g694(.A1(new_n822_), .A2(new_n824_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  AND2_X1   g695(.A1(new_n682_), .A2(G330), .ZN(new_n832_));
  OR2_X1    g696(.A1(new_n648_), .A2(new_n832_), .ZN(new_n833_));
  AOI211_X1 g697(.A(new_n506_), .B(new_n614_), .C1(new_n513_), .C2(new_n521_), .ZN(new_n834_));
  OAI21_X1  g698(.A(new_n654_), .B1(new_n659_), .B2(KEYINPUT45), .ZN(new_n835_));
  OAI211_X1 g699(.A(new_n834_), .B(new_n667_), .C1(new_n825_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g700(.A1(new_n825_), .A2(new_n667_), .ZN(new_n837_));
  NAND2_X1  g701(.A1(new_n513_), .A2(new_n521_), .ZN(new_n838_));
  NAND4_X1  g702(.A1(new_n838_), .A2(G330), .A3(new_n613_), .A4(new_n667_), .ZN(new_n839_));
  INV_X1    g703(.A(new_n835_), .ZN(new_n840_));
  NAND3_X1  g704(.A1(new_n837_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g705(.A1(new_n653_), .A2(KEYINPUT44), .ZN(new_n842_));
  NAND2_X1  g706(.A1(new_n842_), .A2(KEYINPUT45), .ZN(new_n843_));
  INV_X1    g707(.A(new_n843_), .ZN(new_n844_));
  AND3_X1   g708(.A1(new_n836_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g709(.A(new_n844_), .B1(new_n836_), .B2(new_n841_), .ZN(new_n846_));
  OAI22_X1  g710(.A1(new_n831_), .A2(new_n833_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g711(.A1(new_n829_), .A2(KEYINPUT46), .ZN(new_n848_));
  NAND4_X1  g712(.A1(new_n824_), .A2(new_n848_), .A3(new_n834_), .A4(new_n818_), .ZN(new_n849_));
  NAND2_X1  g713(.A1(new_n828_), .A2(new_n830_), .ZN(new_n850_));
  NAND2_X1  g714(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AND3_X1   g715(.A1(new_n837_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n852_));
  AOI21_X1  g716(.A(new_n839_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n853_));
  OAI21_X1  g717(.A(new_n843_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g718(.A1(new_n836_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n855_));
  NOR2_X1   g719(.A1(new_n648_), .A2(new_n832_), .ZN(new_n856_));
  NAND4_X1  g720(.A1(new_n851_), .A2(new_n854_), .A3(new_n855_), .A4(new_n856_), .ZN(new_n857_));
  NAND3_X1  g721(.A1(new_n847_), .A2(new_n857_), .A3(new_n502_), .ZN(new_n858_));
  OAI21_X1  g722(.A(new_n534_), .B1(new_n620_), .B2(G58), .ZN(new_n859_));
  NAND2_X1  g723(.A1(new_n653_), .A2(new_n543_), .ZN(new_n860_));
  XOR2_X1   g724(.A(new_n860_), .B(KEYINPUT49), .Z(new_n861_));
  AOI211_X1 g725(.A(new_n188_), .B(new_n566_), .C1(new_n626_), .C2(G107), .ZN(new_n862_));
  OAI221_X1 g726(.A(new_n862_), .B1(new_n686_), .B2(new_n555_), .C1(new_n582_), .C2(new_n571_), .ZN(new_n863_));
  AOI22_X1  g727(.A1(G283), .A2(new_n795_), .B1(new_n623_), .B2(G97), .ZN(new_n864_));
  OAI221_X1 g728(.A(new_n864_), .B1(new_n138_), .B2(new_n568_), .C1(new_n377_), .C2(new_n562_), .ZN(new_n865_));
  AOI22_X1  g729(.A1(new_n765_), .A2(G132), .B1(G125), .B2(new_n572_), .ZN(new_n866_));
  OAI21_X1  g730(.A(KEYINPUT48), .B1(new_n568_), .B2(new_n203_), .ZN(new_n867_));
  OAI211_X1 g731(.A(new_n866_), .B(new_n867_), .C1(new_n637_), .C2(new_n569_), .ZN(new_n868_));
  AOI21_X1  g732(.A(G33), .B1(new_n623_), .B2(G143), .ZN(new_n869_));
  AOI22_X1  g733(.A1(new_n797_), .A2(G150), .B1(new_n628_), .B2(G159), .ZN(new_n870_));
  NAND2_X1  g734(.A1(new_n795_), .A2(G128), .ZN(new_n871_));
  OR3_X1    g735(.A1(new_n568_), .A2(KEYINPUT48), .A3(new_n203_), .ZN(new_n872_));
  NAND4_X1  g736(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  OAI22_X1  g737(.A1(new_n863_), .A2(new_n865_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n874_));
  AOI211_X1 g738(.A(new_n859_), .B(new_n861_), .C1(new_n546_), .C2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g739(.A1(new_n845_), .A2(new_n846_), .ZN(new_n876_));
  AOI21_X1  g740(.A(new_n875_), .B1(new_n876_), .B2(new_n533_), .ZN(new_n877_));
  NAND2_X1  g741(.A1(new_n858_), .A2(new_n877_), .ZN(G378));
  OAI21_X1  g742(.A(new_n534_), .B1(new_n620_), .B2(G50), .ZN(new_n879_));
  AOI22_X1  g743(.A1(new_n765_), .A2(G107), .B1(G283), .B2(new_n572_), .ZN(new_n880_));
  AOI211_X1 g744(.A(new_n188_), .B(G41), .C1(new_n628_), .C2(G68), .ZN(new_n881_));
  OAI211_X1 g745(.A(new_n880_), .B(new_n881_), .C1(new_n286_), .C2(new_n569_), .ZN(new_n882_));
  NOR2_X1   g746(.A1(new_n568_), .A2(new_n137_), .ZN(new_n883_));
  OAI22_X1  g747(.A1(new_n557_), .A2(new_n686_), .B1(new_n560_), .B2(new_n406_), .ZN(new_n884_));
  NOR4_X1   g748(.A1(new_n882_), .A2(new_n776_), .A3(new_n883_), .A4(new_n884_), .ZN(new_n885_));
  XOR2_X1   g749(.A(new_n885_), .B(KEYINPUT53), .Z(new_n886_));
  INV_X1    g750(.A(G125), .ZN(new_n887_));
  OAI211_X1 g751(.A(new_n188_), .B(new_n173_), .C1(new_n557_), .C2(new_n887_), .ZN(new_n888_));
  INV_X1    g752(.A(G128), .ZN(new_n889_));
  NOR2_X1   g753(.A1(new_n555_), .A2(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g754(.A(KEYINPUT54), .B(G132), .ZN(new_n891_));
  AOI211_X1 g755(.A(new_n888_), .B(new_n890_), .C1(new_n626_), .C2(new_n891_), .ZN(new_n892_));
  INV_X1    g756(.A(KEYINPUT55), .ZN(new_n893_));
  AND3_X1   g757(.A1(new_n572_), .A2(new_n893_), .A3(G124), .ZN(new_n894_));
  AOI21_X1  g758(.A(new_n893_), .B1(new_n572_), .B2(G124), .ZN(new_n895_));
  OAI22_X1  g759(.A1(new_n560_), .A2(new_n637_), .B1(new_n634_), .B2(new_n562_), .ZN(new_n896_));
  OAI22_X1  g760(.A1(new_n633_), .A2(new_n565_), .B1(new_n568_), .B2(new_n733_), .ZN(new_n897_));
  NOR4_X1   g761(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .A4(new_n897_), .ZN(new_n898_));
  AOI22_X1  g762(.A1(new_n892_), .A2(new_n898_), .B1(G41), .B2(new_n203_), .ZN(new_n899_));
  NAND2_X1  g763(.A1(new_n886_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g764(.A(new_n879_), .B1(new_n900_), .B2(new_n546_), .ZN(new_n901_));
  NAND2_X1  g765(.A1(new_n212_), .A2(new_n649_), .ZN(new_n902_));
  XNOR2_X1  g766(.A(new_n226_), .B(new_n902_), .ZN(new_n903_));
  INV_X1    g767(.A(new_n903_), .ZN(new_n904_));
  OR2_X1    g768(.A1(new_n904_), .A2(new_n544_), .ZN(new_n905_));
  NAND2_X1  g769(.A1(new_n901_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g770(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g771(.A1(new_n673_), .A2(new_n675_), .ZN(new_n908_));
  INV_X1    g772(.A(new_n670_), .ZN(new_n909_));
  NAND2_X1  g773(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g774(.A1(new_n910_), .A2(new_n903_), .ZN(new_n911_));
  NAND2_X1  g775(.A1(new_n676_), .A2(new_n904_), .ZN(new_n912_));
  NAND2_X1  g776(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NOR3_X1   g777(.A1(new_n454_), .A2(new_n348_), .A3(new_n483_), .ZN(new_n914_));
  OAI211_X1 g778(.A(new_n681_), .B(G330), .C1(new_n914_), .C2(new_n520_), .ZN(new_n915_));
  INV_X1    g779(.A(KEYINPUT51), .ZN(new_n916_));
  NAND2_X1  g780(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g781(.A1(new_n522_), .A2(KEYINPUT51), .A3(new_n681_), .ZN(new_n918_));
  NAND2_X1  g782(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g783(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g784(.A1(new_n913_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g785(.A1(new_n672_), .A2(new_n671_), .ZN(new_n922_));
  NAND2_X1  g786(.A1(new_n669_), .A2(KEYINPUT50), .ZN(new_n923_));
  INV_X1    g787(.A(KEYINPUT50), .ZN(new_n924_));
  NAND4_X1  g788(.A1(new_n659_), .A2(new_n667_), .A3(new_n924_), .A4(new_n668_), .ZN(new_n925_));
  NAND4_X1  g789(.A1(new_n923_), .A2(new_n656_), .A3(new_n904_), .A4(new_n925_), .ZN(new_n926_));
  OR2_X1    g790(.A1(new_n922_), .A2(new_n926_), .ZN(new_n927_));
  OAI211_X1 g791(.A(new_n919_), .B(new_n927_), .C1(new_n676_), .C2(new_n904_), .ZN(new_n928_));
  INV_X1    g792(.A(KEYINPUT52), .ZN(new_n929_));
  AND2_X1   g793(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g794(.A1(new_n928_), .A2(new_n929_), .ZN(new_n931_));
  OAI21_X1  g795(.A(new_n921_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  AOI21_X1  g796(.A(new_n907_), .B1(new_n932_), .B2(new_n533_), .ZN(new_n933_));
  NAND2_X1  g797(.A1(new_n857_), .A2(new_n856_), .ZN(new_n934_));
  NOR2_X1   g798(.A1(new_n676_), .A2(new_n904_), .ZN(new_n935_));
  INV_X1    g799(.A(new_n927_), .ZN(new_n936_));
  OAI21_X1  g800(.A(new_n920_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g801(.A1(new_n937_), .A2(new_n928_), .ZN(new_n938_));
  NAND3_X1  g802(.A1(new_n934_), .A2(new_n502_), .A3(new_n938_), .ZN(new_n939_));
  NAND2_X1  g803(.A1(new_n933_), .A2(new_n939_), .ZN(G375));
  NAND2_X1  g804(.A1(new_n671_), .A2(new_n543_), .ZN(new_n941_));
  OAI21_X1  g805(.A(new_n534_), .B1(new_n620_), .B2(G68), .ZN(new_n942_));
  AOI211_X1 g806(.A(G33), .B(new_n883_), .C1(new_n626_), .C2(G143), .ZN(new_n943_));
  OAI221_X1 g807(.A(new_n943_), .B1(new_n889_), .B2(new_n571_), .C1(new_n637_), .C2(new_n555_), .ZN(new_n944_));
  AOI22_X1  g808(.A1(new_n795_), .A2(G132), .B1(new_n628_), .B2(G50), .ZN(new_n945_));
  OAI221_X1 g809(.A(new_n945_), .B1(new_n634_), .B2(new_n560_), .C1(new_n733_), .C2(new_n565_), .ZN(new_n946_));
  AOI21_X1  g810(.A(new_n775_), .B1(new_n623_), .B2(G107), .ZN(new_n947_));
  OAI221_X1 g811(.A(new_n947_), .B1(new_n286_), .B2(new_n565_), .C1(new_n582_), .C2(new_n557_), .ZN(new_n948_));
  OAI21_X1  g812(.A(G33), .B1(new_n568_), .B2(new_n377_), .ZN(new_n949_));
  AOI21_X1  g813(.A(new_n949_), .B1(new_n626_), .B2(G116), .ZN(new_n950_));
  OAI221_X1 g814(.A(new_n950_), .B1(new_n575_), .B2(new_n555_), .C1(new_n314_), .C2(new_n571_), .ZN(new_n951_));
  OAI22_X1  g815(.A1(new_n944_), .A2(new_n946_), .B1(new_n948_), .B2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g816(.A(new_n942_), .B1(new_n952_), .B2(new_n546_), .ZN(new_n953_));
  AOI22_X1  g817(.A1(new_n851_), .A2(new_n533_), .B1(new_n941_), .B2(new_n953_), .ZN(new_n954_));
  OAI21_X1  g818(.A(new_n502_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n955_));
  NOR2_X1   g819(.A1(new_n851_), .A2(new_n856_), .ZN(new_n956_));
  OAI21_X1  g820(.A(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(G381));
  OR3_X1    g821(.A1(G378), .A2(G384), .A3(G381), .ZN(new_n958_));
  INV_X1    g822(.A(KEYINPUT56), .ZN(new_n959_));
  OR3_X1    g823(.A1(new_n958_), .A2(new_n959_), .A3(G375), .ZN(new_n960_));
  OAI21_X1  g824(.A(new_n959_), .B1(new_n958_), .B2(G375), .ZN(new_n961_));
  NAND2_X1  g825(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  NAND3_X1  g826(.A1(new_n815_), .A2(new_n727_), .A3(new_n749_), .ZN(new_n963_));
  NOR3_X1   g827(.A1(new_n963_), .A2(G396), .A3(G393), .ZN(new_n964_));
  AND3_X1   g828(.A1(new_n962_), .A2(KEYINPUT57), .A3(new_n964_), .ZN(new_n965_));
  AOI21_X1  g829(.A(KEYINPUT57), .B1(new_n962_), .B2(new_n964_), .ZN(new_n966_));
  OR2_X1    g830(.A1(new_n965_), .A2(new_n966_), .ZN(G407));
  AOI221_X4 g831(.A(new_n503_), .B1(new_n928_), .B2(new_n937_), .C1(new_n857_), .C2(new_n856_), .ZN(new_n968_));
  NAND4_X1  g832(.A1(new_n911_), .A2(KEYINPUT52), .A3(new_n919_), .A4(new_n927_), .ZN(new_n969_));
  NAND2_X1  g833(.A1(new_n928_), .A2(new_n929_), .ZN(new_n970_));
  AOI22_X1  g834(.A1(new_n969_), .A2(new_n970_), .B1(new_n913_), .B2(new_n920_), .ZN(new_n971_));
  OAI21_X1  g835(.A(new_n906_), .B1(new_n971_), .B2(new_n532_), .ZN(new_n972_));
  NOR2_X1   g836(.A1(new_n968_), .A2(new_n972_), .ZN(new_n973_));
  NAND4_X1  g837(.A1(new_n973_), .A2(new_n482_), .A3(new_n858_), .A4(new_n877_), .ZN(new_n974_));
  OAI211_X1 g838(.A(G213), .B(new_n974_), .C1(new_n965_), .C2(new_n966_), .ZN(G409));
  NAND2_X1  g839(.A1(new_n482_), .A2(G213), .ZN(new_n976_));
  NAND3_X1  g840(.A1(new_n858_), .A2(new_n877_), .A3(new_n976_), .ZN(new_n977_));
  NOR2_X1   g841(.A1(new_n971_), .A2(new_n857_), .ZN(new_n978_));
  AOI21_X1  g842(.A(new_n856_), .B1(new_n937_), .B2(new_n928_), .ZN(new_n979_));
  OAI21_X1  g843(.A(new_n502_), .B1(new_n978_), .B2(new_n979_), .ZN(new_n980_));
  AOI21_X1  g844(.A(new_n977_), .B1(new_n980_), .B2(new_n933_), .ZN(new_n981_));
  NAND4_X1  g845(.A1(new_n973_), .A2(KEYINPUT58), .A3(G378), .A4(new_n976_), .ZN(new_n982_));
  NAND4_X1  g846(.A1(new_n933_), .A2(G378), .A3(new_n939_), .A4(new_n976_), .ZN(new_n983_));
  INV_X1    g847(.A(KEYINPUT58), .ZN(new_n984_));
  NAND2_X1  g848(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  AOI21_X1  g849(.A(new_n981_), .B1(new_n982_), .B2(new_n985_), .ZN(new_n986_));
  INV_X1    g850(.A(KEYINPUT61), .ZN(new_n987_));
  INV_X1    g851(.A(KEYINPUT59), .ZN(new_n988_));
  OAI21_X1  g852(.A(new_n988_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n989_));
  AOI21_X1  g853(.A(new_n503_), .B1(new_n851_), .B2(new_n856_), .ZN(new_n990_));
  NAND2_X1  g854(.A1(new_n831_), .A2(new_n833_), .ZN(new_n991_));
  NAND3_X1  g855(.A1(new_n990_), .A2(KEYINPUT59), .A3(new_n991_), .ZN(new_n992_));
  NAND2_X1  g856(.A1(new_n989_), .A2(new_n992_), .ZN(new_n993_));
  AOI21_X1  g857(.A(G384), .B1(new_n993_), .B2(new_n954_), .ZN(new_n994_));
  INV_X1    g858(.A(new_n954_), .ZN(new_n995_));
  AOI211_X1 g859(.A(new_n644_), .B(new_n995_), .C1(new_n989_), .C2(new_n992_), .ZN(new_n996_));
  NOR2_X1   g860(.A1(new_n994_), .A2(new_n996_), .ZN(new_n997_));
  NAND3_X1  g861(.A1(new_n482_), .A2(G213), .A3(G2897), .ZN(new_n998_));
  INV_X1    g862(.A(new_n998_), .ZN(new_n999_));
  AOI21_X1  g863(.A(new_n987_), .B1(new_n997_), .B2(new_n999_), .ZN(new_n1000_));
  NOR4_X1   g864(.A1(new_n994_), .A2(new_n996_), .A3(KEYINPUT61), .A4(new_n998_), .ZN(new_n1001_));
  OAI21_X1  g865(.A(new_n986_), .B1(new_n1000_), .B2(new_n1001_), .ZN(new_n1002_));
  NAND2_X1  g866(.A1(new_n980_), .A2(new_n933_), .ZN(new_n1003_));
  INV_X1    g867(.A(new_n977_), .ZN(new_n1004_));
  NAND2_X1  g868(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1005_));
  AND2_X1   g869(.A1(new_n983_), .A2(new_n984_), .ZN(new_n1006_));
  NOR2_X1   g870(.A1(new_n983_), .A2(new_n984_), .ZN(new_n1007_));
  OAI21_X1  g871(.A(new_n1005_), .B1(new_n1006_), .B2(new_n1007_), .ZN(new_n1008_));
  INV_X1    g872(.A(KEYINPUT60), .ZN(new_n1009_));
  AOI21_X1  g873(.A(new_n995_), .B1(new_n989_), .B2(new_n992_), .ZN(new_n1010_));
  AOI21_X1  g874(.A(new_n1009_), .B1(new_n1010_), .B2(G384), .ZN(new_n1011_));
  OAI22_X1  g875(.A1(new_n1011_), .A2(new_n999_), .B1(new_n994_), .B2(new_n996_), .ZN(new_n1012_));
  INV_X1    g876(.A(new_n992_), .ZN(new_n1013_));
  AOI21_X1  g877(.A(KEYINPUT59), .B1(new_n990_), .B2(new_n991_), .ZN(new_n1014_));
  OAI21_X1  g878(.A(new_n954_), .B1(new_n1013_), .B2(new_n1014_), .ZN(new_n1015_));
  NAND2_X1  g879(.A1(new_n1015_), .A2(new_n644_), .ZN(new_n1016_));
  NAND2_X1  g880(.A1(new_n1010_), .A2(G384), .ZN(new_n1017_));
  NAND4_X1  g881(.A1(new_n1016_), .A2(new_n1017_), .A3(new_n1009_), .A4(new_n998_), .ZN(new_n1018_));
  NAND2_X1  g882(.A1(new_n1012_), .A2(new_n1018_), .ZN(new_n1019_));
  NAND2_X1  g883(.A1(new_n1008_), .A2(new_n1019_), .ZN(new_n1020_));
  INV_X1    g884(.A(new_n997_), .ZN(new_n1021_));
  NAND3_X1  g885(.A1(new_n986_), .A2(new_n1021_), .A3(new_n998_), .ZN(new_n1022_));
  NAND3_X1  g886(.A1(new_n1002_), .A2(new_n1020_), .A3(new_n1022_), .ZN(new_n1023_));
  AND2_X1   g887(.A1(G393), .A2(G396), .ZN(new_n1024_));
  NOR2_X1   g888(.A1(G393), .A2(G396), .ZN(new_n1025_));
  NOR2_X1   g889(.A1(new_n1024_), .A2(new_n1025_), .ZN(new_n1026_));
  AND3_X1   g890(.A1(new_n815_), .A2(new_n727_), .A3(new_n749_), .ZN(new_n1027_));
  NAND2_X1  g891(.A1(new_n810_), .A2(new_n814_), .ZN(new_n1028_));
  NAND2_X1  g892(.A1(new_n787_), .A2(new_n789_), .ZN(new_n1029_));
  AOI22_X1  g893(.A1(new_n727_), .A2(new_n749_), .B1(new_n1028_), .B2(new_n1029_), .ZN(new_n1030_));
  OAI21_X1  g894(.A(new_n1026_), .B1(new_n1027_), .B2(new_n1030_), .ZN(new_n1031_));
  NAND2_X1  g895(.A1(G390), .A2(G387), .ZN(new_n1032_));
  OR2_X1    g896(.A1(new_n1024_), .A2(new_n1025_), .ZN(new_n1033_));
  NAND3_X1  g897(.A1(new_n1032_), .A2(new_n1033_), .A3(new_n963_), .ZN(new_n1034_));
  INV_X1    g898(.A(KEYINPUT62), .ZN(new_n1035_));
  NAND3_X1  g899(.A1(new_n1031_), .A2(new_n1034_), .A3(new_n1035_), .ZN(new_n1036_));
  NAND4_X1  g900(.A1(new_n1032_), .A2(new_n1033_), .A3(KEYINPUT62), .A4(new_n963_), .ZN(new_n1037_));
  NAND2_X1  g901(.A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1038_));
  INV_X1    g902(.A(new_n1038_), .ZN(new_n1039_));
  NAND2_X1  g903(.A1(new_n1023_), .A2(new_n1039_), .ZN(new_n1040_));
  NAND2_X1  g904(.A1(new_n1002_), .A2(KEYINPUT63), .ZN(new_n1041_));
  INV_X1    g905(.A(KEYINPUT63), .ZN(new_n1042_));
  OAI211_X1 g906(.A(new_n986_), .B(new_n1042_), .C1(new_n1000_), .C2(new_n1001_), .ZN(new_n1043_));
  NAND2_X1  g907(.A1(new_n1041_), .A2(new_n1043_), .ZN(new_n1044_));
  NAND4_X1  g908(.A1(new_n1020_), .A2(new_n1022_), .A3(new_n1034_), .A4(new_n1031_), .ZN(new_n1045_));
  OAI21_X1  g909(.A(new_n1040_), .B1(new_n1044_), .B2(new_n1045_), .ZN(G405));
  XNOR2_X1  g910(.A(new_n973_), .B(G378), .ZN(new_n1047_));
  NAND3_X1  g911(.A1(new_n1036_), .A2(new_n1037_), .A3(new_n1047_), .ZN(new_n1048_));
  INV_X1    g912(.A(new_n1048_), .ZN(new_n1049_));
  AOI21_X1  g913(.A(new_n1047_), .B1(new_n1036_), .B2(new_n1037_), .ZN(new_n1050_));
  NOR3_X1   g914(.A1(new_n1049_), .A2(new_n1050_), .A3(new_n1021_), .ZN(new_n1051_));
  INV_X1    g915(.A(new_n1047_), .ZN(new_n1052_));
  NAND2_X1  g916(.A1(new_n1038_), .A2(new_n1052_), .ZN(new_n1053_));
  AOI21_X1  g917(.A(new_n997_), .B1(new_n1053_), .B2(new_n1048_), .ZN(new_n1054_));
  NOR2_X1   g918(.A1(new_n1051_), .A2(new_n1054_), .ZN(G402));
endmodule


