//Secret key is'0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_c5315" written by ABC on Wed Nov 16 10:39:49 2022

module locked_c5315 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G4, G11, G14, G17, G20, G23, G24, G25,
    G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64,
    G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94,
    G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161,
    G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197,
    G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241,
    G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281,
    G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324,
    G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372,
    G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479,
    G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562,
    G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546,
    G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091,
    G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G4, G11, G14, G17, G20, G23,
    G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54,
    G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88,
    G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116,
    G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130,
    G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155,
    G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191,
    G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233,
    G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273,
    G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316,
    G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366,
    G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457,
    G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559,
    G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173,
    G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090,
    G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_n444_, new_n449_, new_n451_, new_n461_, new_n469_, new_n470_,
    new_n472_, new_n476_, new_n477_, new_n478_, new_n480_, new_n481_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n490_, new_n491_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1104_, new_n1105_,
    new_n1106_, new_n1108_, new_n1109_, new_n1110_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1118_, new_n1119_, new_n1120_,
    new_n1122_, new_n1123_, new_n1124_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1198_, new_n1199_,
    new_n1201_, new_n1202_, new_n1203_, new_n1205_, new_n1206_, new_n1207_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1215_,
    new_n1216_, new_n1218_, new_n1219_, new_n1220_, new_n1222_, new_n1223_,
    new_n1224_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1244_, new_n1245_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1263_, new_n1264_, new_n1265_, new_n1267_, new_n1268_,
    new_n1269_, new_n1271_, new_n1272_, new_n1273_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_;
  BUF_X1    g0000(.A(G141), .Z(G144));
  BUF_X1    g0001(.A(G293), .Z(G298));
  BUF_X1    g0002(.A(G3173), .Z(G973));
  INV_X1    g0003(.A(G545), .ZN(G594));
  INV_X1    g0004(.A(G348), .ZN(G599));
  INV_X1    g0005(.A(G366), .ZN(G600));
  INV_X1    g0006(.A(G552), .ZN(G849));
  INV_X1    g0007(.A(G562), .ZN(G850));
  NOR2_X1   g0008(.A1(G849), .A2(G850), .ZN(G601));
  INV_X1    g0009(.A(G549), .ZN(G602));
  INV_X1    g0010(.A(G545), .ZN(G603));
  INV_X1    g0011(.A(G545), .ZN(G604));
  XNOR2_X1  g0012(.A(KEYINPUT0), .B(G338), .ZN(G611));
  INV_X1    g0013(.A(G358), .ZN(G612));
  NAND2_X1  g0014(.A1(G141), .A2(G145), .ZN(new_n444_));
  XNOR2_X1  g0015(.A(new_n444_), .B(KEYINPUT1), .ZN(G810));
  INV_X1    g0016(.A(G245), .ZN(G848));
  INV_X1    g0017(.A(G559), .ZN(G851));
  AND2_X1   g0018(.A1(G1), .A2(G373), .ZN(G634));
  INV_X1    g0019(.A(G136), .ZN(new_n449_));
  NOR2_X1   g0020(.A1(new_n449_), .A2(G3173), .ZN(G815));
  INV_X1    g0021(.A(G2824), .ZN(new_n451_));
  NAND2_X1  g0022(.A1(new_n451_), .A2(G27), .ZN(G845));
  NAND2_X1  g0023(.A1(G386), .A2(G556), .ZN(G847));
  BUF_X1    g0024(.A(G137), .Z(G926));
  BUF_X1    g0025(.A(G141), .Z(G923));
  BUF_X1    g0026(.A(G1), .Z(G921));
  BUF_X1    g0027(.A(G549), .Z(G892));
  BUF_X1    g0028(.A(G299), .Z(G887));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G549), .Z(G606));
  NAND2_X1  g0030(.A1(G27), .A2(G31), .ZN(G809));
  INV_X1    g0031(.A(G809), .ZN(new_n461_));
  NAND2_X1  g0032(.A1(new_n461_), .A2(G140), .ZN(G656));
  XNOR2_X1  g0033(.A(KEYINPUT3), .B(G1), .ZN(G993));
  BUF_X1    g0034(.A(G1), .Z(G978));
  BUF_X1    g0035(.A(G1), .Z(G949));
  XNOR2_X1  g0036(.A(KEYINPUT4), .B(G1), .ZN(G939));
  BUF_X1    g0037(.A(G299), .Z(G889));
  INV_X1    g0038(.A(G299), .ZN(G593));
  OR2_X1    g0039(.A1(G86), .A2(G2358), .ZN(new_n469_));
  INV_X1    g0040(.A(G2358), .ZN(new_n470_));
  OAI211_X1 g0041(.A(new_n469_), .B(new_n461_), .C1(G87), .C2(new_n470_), .ZN(G636));
  OR2_X1    g0042(.A1(G88), .A2(G2358), .ZN(new_n472_));
  OAI211_X1 g0043(.A(new_n472_), .B(new_n461_), .C1(G34), .C2(new_n470_), .ZN(G704));
  OAI211_X1 g0044(.A(new_n472_), .B(new_n461_), .C1(G34), .C2(new_n470_), .ZN(G717));
  NAND2_X1  g0045(.A1(new_n461_), .A2(G83), .ZN(G820));
  INV_X1    g0046(.A(G141), .ZN(new_n476_));
  AOI21_X1  g0047(.A(G809), .B1(G24), .B2(new_n470_), .ZN(new_n477_));
  NAND2_X1  g0048(.A1(G25), .A2(G2358), .ZN(new_n478_));
  AOI21_X1  g0049(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(G639));
  AOI21_X1  g0050(.A(G809), .B1(G26), .B2(new_n470_), .ZN(new_n480_));
  NAND2_X1  g0051(.A1(G81), .A2(G2358), .ZN(new_n481_));
  AOI21_X1  g0052(.A(new_n476_), .B1(new_n480_), .B2(new_n481_), .ZN(G673));
  INV_X1    g0053(.A(G79), .ZN(new_n483_));
  OAI21_X1  g0054(.A(new_n461_), .B1(new_n483_), .B2(G2358), .ZN(new_n484_));
  INV_X1    g0055(.A(KEYINPUT5), .ZN(new_n485_));
  OR2_X1    g0056(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AND2_X1   g0057(.A1(G23), .A2(G2358), .ZN(new_n487_));
  AOI22_X1  g0058(.A1(new_n484_), .A2(new_n485_), .B1(new_n461_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g0059(.A(new_n476_), .B1(new_n486_), .B2(new_n488_), .ZN(G707));
  AOI21_X1  g0060(.A(G809), .B1(G82), .B2(new_n470_), .ZN(new_n490_));
  NAND2_X1  g0061(.A1(G80), .A2(G2358), .ZN(new_n491_));
  AOI21_X1  g0062(.A(new_n476_), .B1(new_n490_), .B2(new_n491_), .ZN(G715));
  INV_X1    g0063(.A(G3552), .ZN(new_n493_));
  OR2_X1    g0064(.A1(new_n493_), .A2(KEYINPUT6), .ZN(new_n494_));
  NAND2_X1  g0065(.A1(new_n493_), .A2(KEYINPUT6), .ZN(new_n495_));
  NAND2_X1  g0066(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g0067(.A(G351), .ZN(new_n497_));
  OAI21_X1  g0068(.A(G534), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g0069(.A(G3550), .ZN(new_n499_));
  XNOR2_X1  g0070(.A(KEYINPUT7), .B(G351), .ZN(new_n500_));
  AOI21_X1  g0071(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g0072(.A(G534), .ZN(new_n502_));
  OAI22_X1  g0073(.A1(new_n500_), .A2(G3546), .B1(G351), .B2(G3548), .ZN(new_n503_));
  AOI21_X1  g0074(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g0075(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g0076(.A(G523), .B1(G341), .B2(G3550), .ZN(new_n506_));
  INV_X1    g0077(.A(new_n496_), .ZN(new_n507_));
  AOI21_X1  g0078(.A(new_n506_), .B1(new_n507_), .B2(G341), .ZN(new_n508_));
  NAND2_X1  g0079(.A1(G341), .A2(G3546), .ZN(new_n509_));
  INV_X1    g0080(.A(G341), .ZN(new_n510_));
  AOI21_X1  g0081(.A(G523), .B1(new_n510_), .B2(G3548), .ZN(new_n511_));
  AOI21_X1  g0082(.A(new_n508_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g0083(.A1(G254), .A2(G293), .ZN(new_n513_));
  INV_X1    g0084(.A(G242), .ZN(new_n514_));
  AOI21_X1  g0085(.A(new_n513_), .B1(new_n514_), .B2(G293), .ZN(new_n515_));
  INV_X1    g0086(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g0087(.A1(G251), .A2(G302), .ZN(new_n517_));
  INV_X1    g0088(.A(G248), .ZN(new_n518_));
  AOI21_X1  g0089(.A(new_n517_), .B1(new_n518_), .B2(G302), .ZN(new_n519_));
  AND2_X1   g0090(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g0091(.A1(G251), .A2(G361), .ZN(new_n521_));
  AOI21_X1  g0092(.A(new_n521_), .B1(new_n518_), .B2(G361), .ZN(new_n522_));
  NOR2_X1   g0093(.A1(G514), .A2(G3546), .ZN(new_n523_));
  AOI21_X1  g0094(.A(new_n523_), .B1(G514), .B2(G3552), .ZN(new_n524_));
  NAND4_X1  g0095(.A1(new_n512_), .A2(new_n520_), .A3(new_n522_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g0096(.A(G324), .ZN(new_n526_));
  NAND3_X1  g0097(.A1(new_n526_), .A2(new_n499_), .A3(G503), .ZN(new_n527_));
  XNOR2_X1  g0098(.A(new_n527_), .B(KEYINPUT8), .ZN(new_n528_));
  INV_X1    g0099(.A(G503), .ZN(new_n529_));
  NOR3_X1   g0100(.A1(new_n496_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g0101(.A(G3546), .ZN(new_n531_));
  NAND2_X1  g0102(.A1(new_n531_), .A2(G324), .ZN(new_n532_));
  INV_X1    g0103(.A(G3548), .ZN(new_n533_));
  AOI21_X1  g0104(.A(G503), .B1(new_n526_), .B2(new_n533_), .ZN(new_n534_));
  AOI211_X1 g0105(.A(new_n528_), .B(new_n530_), .C1(new_n532_), .C2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g0106(.A1(G248), .A2(G308), .ZN(new_n536_));
  INV_X1    g0107(.A(G479), .ZN(new_n537_));
  INV_X1    g0108(.A(G308), .ZN(new_n538_));
  AOI21_X1  g0109(.A(new_n537_), .B1(G251), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g0110(.A(G254), .ZN(new_n540_));
  AOI21_X1  g0111(.A(G479), .B1(new_n540_), .B2(new_n538_), .ZN(new_n541_));
  NAND2_X1  g0112(.A1(new_n514_), .A2(G308), .ZN(new_n542_));
  AOI22_X1  g0113(.A1(new_n536_), .A2(new_n539_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g0114(.A1(G248), .A2(G316), .ZN(new_n544_));
  INV_X1    g0115(.A(G251), .ZN(new_n545_));
  OAI211_X1 g0116(.A(new_n544_), .B(G490), .C1(new_n545_), .C2(G316), .ZN(new_n546_));
  INV_X1    g0117(.A(G316), .ZN(new_n547_));
  AOI21_X1  g0118(.A(G490), .B1(new_n540_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g0119(.A(new_n548_), .B1(G242), .B2(new_n547_), .ZN(new_n549_));
  NAND3_X1  g0120(.A1(new_n543_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  NOR4_X1   g0121(.A1(new_n505_), .A2(new_n525_), .A3(new_n535_), .A4(new_n550_), .ZN(G598));
  OAI21_X1  g0122(.A(G400), .B1(G265), .B2(G3550), .ZN(new_n552_));
  AOI21_X1  g0123(.A(new_n552_), .B1(new_n507_), .B2(G265), .ZN(new_n553_));
  NAND2_X1  g0124(.A1(G265), .A2(G3546), .ZN(new_n554_));
  INV_X1    g0125(.A(G265), .ZN(new_n555_));
  AOI21_X1  g0126(.A(G400), .B1(new_n555_), .B2(G3548), .ZN(new_n556_));
  AOI21_X1  g0127(.A(new_n553_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g0128(.A(G374), .ZN(new_n558_));
  INV_X1    g0129(.A(G281), .ZN(new_n559_));
  OAI21_X1  g0130(.A(new_n558_), .B1(new_n559_), .B2(G3546), .ZN(new_n560_));
  INV_X1    g0131(.A(KEYINPUT13), .ZN(new_n561_));
  OAI22_X1  g0132(.A1(new_n560_), .A2(new_n561_), .B1(G281), .B2(G3548), .ZN(new_n562_));
  AOI21_X1  g0133(.A(new_n562_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n563_));
  OAI21_X1  g0134(.A(G374), .B1(new_n499_), .B2(G281), .ZN(new_n564_));
  AOI21_X1  g0135(.A(new_n564_), .B1(new_n496_), .B2(G281), .ZN(new_n565_));
  OR2_X1    g0136(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g0137(.A(G389), .ZN(new_n567_));
  INV_X1    g0138(.A(G257), .ZN(new_n568_));
  AOI21_X1  g0139(.A(new_n567_), .B1(new_n568_), .B2(G3550), .ZN(new_n569_));
  OAI21_X1  g0140(.A(new_n569_), .B1(new_n507_), .B2(new_n568_), .ZN(new_n570_));
  OAI21_X1  g0141(.A(new_n567_), .B1(new_n568_), .B2(G3546), .ZN(new_n571_));
  AOI22_X1  g0142(.A1(new_n571_), .A2(KEYINPUT14), .B1(new_n568_), .B2(new_n533_), .ZN(new_n572_));
  OAI21_X1  g0143(.A(new_n572_), .B1(KEYINPUT14), .B2(new_n571_), .ZN(new_n573_));
  NAND2_X1  g0144(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g0145(.A(G411), .B1(G273), .B2(G3550), .ZN(new_n575_));
  AOI21_X1  g0146(.A(new_n575_), .B1(new_n507_), .B2(G273), .ZN(new_n576_));
  INV_X1    g0147(.A(G411), .ZN(new_n577_));
  OAI21_X1  g0148(.A(new_n577_), .B1(new_n533_), .B2(G273), .ZN(new_n578_));
  AOI21_X1  g0149(.A(new_n578_), .B1(G273), .B2(G3546), .ZN(new_n579_));
  NOR2_X1   g0150(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g0151(.A1(new_n557_), .A2(new_n566_), .A3(new_n574_), .A4(new_n580_), .ZN(new_n581_));
  OR2_X1    g0152(.A1(new_n581_), .A2(KEYINPUT15), .ZN(new_n582_));
  NAND3_X1  g0153(.A1(G206), .A2(G248), .A3(G446), .ZN(new_n583_));
  XOR2_X1   g0154(.A(new_n583_), .B(KEYINPUT16), .Z(new_n584_));
  INV_X1    g0155(.A(G446), .ZN(new_n585_));
  NOR3_X1   g0156(.A1(new_n545_), .A2(new_n585_), .A3(G206), .ZN(new_n586_));
  OAI21_X1  g0157(.A(new_n585_), .B1(new_n540_), .B2(G206), .ZN(new_n587_));
  AOI21_X1  g0158(.A(new_n587_), .B1(G206), .B2(G242), .ZN(new_n588_));
  OR3_X1    g0159(.A1(new_n584_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  XOR2_X1   g0160(.A(new_n589_), .B(KEYINPUT17), .Z(new_n590_));
  INV_X1    g0161(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g0162(.A(G435), .ZN(new_n592_));
  OR2_X1    g0163(.A1(new_n592_), .A2(G234), .ZN(new_n593_));
  OR2_X1    g0164(.A1(new_n593_), .A2(G3550), .ZN(new_n594_));
  NAND2_X1  g0165(.A1(G234), .A2(G435), .ZN(new_n595_));
  AOI21_X1  g0166(.A(G435), .B1(new_n531_), .B2(G234), .ZN(new_n596_));
  INV_X1    g0167(.A(KEYINPUT10), .ZN(new_n597_));
  OAI22_X1  g0168(.A1(new_n596_), .A2(new_n597_), .B1(G234), .B2(G3548), .ZN(new_n598_));
  AND2_X1   g0169(.A1(new_n596_), .A2(new_n597_), .ZN(new_n599_));
  OAI221_X1 g0170(.A(new_n594_), .B1(new_n496_), .B2(new_n595_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g0171(.A1(new_n531_), .A2(G218), .ZN(new_n601_));
  INV_X1    g0172(.A(G468), .ZN(new_n602_));
  OAI211_X1 g0173(.A(new_n601_), .B(new_n602_), .C1(G218), .C2(G3548), .ZN(new_n603_));
  NAND2_X1  g0174(.A1(G218), .A2(G468), .ZN(new_n604_));
  NOR2_X1   g0175(.A1(new_n602_), .A2(G218), .ZN(new_n605_));
  XNOR2_X1  g0176(.A(new_n605_), .B(KEYINPUT9), .ZN(new_n606_));
  OAI221_X1 g0177(.A(new_n603_), .B1(new_n496_), .B2(new_n604_), .C1(new_n606_), .C2(G3550), .ZN(new_n607_));
  INV_X1    g0178(.A(G226), .ZN(new_n608_));
  AOI21_X1  g0179(.A(G422), .B1(new_n608_), .B2(new_n533_), .ZN(new_n609_));
  OAI21_X1  g0180(.A(new_n609_), .B1(new_n608_), .B2(G3546), .ZN(new_n610_));
  NAND2_X1  g0181(.A1(new_n608_), .A2(G422), .ZN(new_n611_));
  NAND2_X1  g0182(.A1(G226), .A2(G422), .ZN(new_n612_));
  OAI221_X1 g0183(.A(new_n610_), .B1(G3550), .B2(new_n611_), .C1(new_n496_), .C2(new_n612_), .ZN(new_n613_));
  AND4_X1   g0184(.A1(new_n591_), .A2(new_n600_), .A3(new_n607_), .A4(new_n613_), .ZN(new_n614_));
  NAND2_X1  g0185(.A1(new_n581_), .A2(KEYINPUT15), .ZN(new_n615_));
  INV_X1    g0186(.A(G210), .ZN(new_n616_));
  XOR2_X1   g0187(.A(KEYINPUT11), .B(G210), .Z(new_n617_));
  INV_X1    g0188(.A(new_n617_), .ZN(new_n618_));
  OAI221_X1 g0189(.A(G457), .B1(new_n496_), .B2(new_n616_), .C1(new_n618_), .C2(G3550), .ZN(new_n619_));
  INV_X1    g0190(.A(G457), .ZN(new_n620_));
  NOR2_X1   g0191(.A1(new_n617_), .A2(G3546), .ZN(new_n621_));
  NOR2_X1   g0192(.A1(G210), .A2(G3548), .ZN(new_n622_));
  OAI21_X1  g0193(.A(new_n620_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g0194(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g0195(.A(new_n624_), .B(KEYINPUT12), .Z(new_n625_));
  AND4_X1   g0196(.A1(new_n582_), .A2(new_n614_), .A3(new_n615_), .A4(new_n625_), .ZN(G610));
  MUX2_X1   g0197(.A(G234), .B(G241), .S(G335), .Z(new_n627_));
  XOR2_X1   g0198(.A(new_n627_), .B(KEYINPUT21), .Z(new_n628_));
  XNOR2_X1  g0199(.A(new_n628_), .B(G435), .ZN(new_n629_));
  INV_X1    g0200(.A(G335), .ZN(new_n630_));
  NOR2_X1   g0201(.A1(new_n630_), .A2(G264), .ZN(new_n631_));
  NOR2_X1   g0202(.A1(G257), .A2(G335), .ZN(new_n632_));
  NOR3_X1   g0203(.A1(new_n631_), .A2(KEYINPUT18), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n634_));
  NAND2_X1  g0205(.A1(new_n568_), .A2(new_n630_), .ZN(new_n635_));
  INV_X1    g0206(.A(G264), .ZN(new_n636_));
  NAND2_X1  g0207(.A1(new_n636_), .A2(G335), .ZN(new_n637_));
  AOI21_X1  g0208(.A(new_n634_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g0209(.A(new_n567_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g0210(.A(KEYINPUT18), .B1(new_n631_), .B2(new_n632_), .ZN(new_n640_));
  NAND3_X1  g0211(.A1(new_n635_), .A2(new_n637_), .A3(new_n634_), .ZN(new_n641_));
  NAND3_X1  g0212(.A1(new_n640_), .A2(new_n641_), .A3(G389), .ZN(new_n642_));
  NAND2_X1  g0213(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g0214(.A(new_n643_), .B(KEYINPUT19), .ZN(new_n644_));
  NAND2_X1  g0215(.A1(new_n629_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g0216(.A1(G288), .A2(G335), .ZN(new_n646_));
  NAND2_X1  g0217(.A1(new_n630_), .A2(KEYINPUT20), .ZN(new_n647_));
  INV_X1    g0218(.A(KEYINPUT20), .ZN(new_n648_));
  NAND2_X1  g0219(.A1(new_n648_), .A2(G335), .ZN(new_n649_));
  NAND2_X1  g0220(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g0221(.A(new_n646_), .B1(new_n650_), .B2(new_n559_), .ZN(new_n651_));
  INV_X1    g0222(.A(KEYINPUT23), .ZN(new_n652_));
  NOR2_X1   g0223(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g0224(.A(KEYINPUT20), .B(G335), .ZN(new_n654_));
  NAND2_X1  g0225(.A1(new_n654_), .A2(G281), .ZN(new_n655_));
  AOI21_X1  g0226(.A(KEYINPUT23), .B1(new_n655_), .B2(new_n646_), .ZN(new_n656_));
  OAI21_X1  g0227(.A(new_n558_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g0228(.A1(G280), .A2(G335), .ZN(new_n658_));
  INV_X1    g0229(.A(G273), .ZN(new_n659_));
  OAI211_X1 g0230(.A(new_n658_), .B(G411), .C1(new_n659_), .C2(G335), .ZN(new_n660_));
  INV_X1    g0231(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0232(.A1(new_n630_), .A2(G273), .ZN(new_n662_));
  AOI21_X1  g0233(.A(G411), .B1(new_n662_), .B2(new_n658_), .ZN(new_n663_));
  OAI21_X1  g0234(.A(KEYINPUT22), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g0235(.A(new_n658_), .B1(new_n659_), .B2(G335), .ZN(new_n665_));
  NAND2_X1  g0236(.A1(new_n665_), .A2(new_n577_), .ZN(new_n666_));
  INV_X1    g0237(.A(KEYINPUT22), .ZN(new_n667_));
  NAND3_X1  g0238(.A1(new_n666_), .A2(new_n667_), .A3(new_n660_), .ZN(new_n668_));
  NAND2_X1  g0239(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g0240(.A1(new_n651_), .A2(new_n652_), .ZN(new_n670_));
  NAND3_X1  g0241(.A1(new_n655_), .A2(KEYINPUT23), .A3(new_n646_), .ZN(new_n671_));
  NAND3_X1  g0242(.A1(new_n670_), .A2(G374), .A3(new_n671_), .ZN(new_n672_));
  NAND3_X1  g0243(.A1(new_n657_), .A2(new_n669_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g0244(.A(G400), .B1(G272), .B2(G335), .ZN(new_n674_));
  OAI21_X1  g0245(.A(new_n674_), .B1(new_n650_), .B2(new_n555_), .ZN(new_n675_));
  INV_X1    g0246(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g0247(.A1(new_n630_), .A2(G265), .ZN(new_n677_));
  NAND2_X1  g0248(.A1(G272), .A2(G335), .ZN(new_n678_));
  NAND2_X1  g0249(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g0250(.A1(new_n679_), .A2(G400), .ZN(new_n680_));
  INV_X1    g0251(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g0252(.A1(new_n676_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g0253(.A(new_n682_), .ZN(new_n683_));
  NOR3_X1   g0254(.A1(new_n645_), .A2(new_n673_), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g0255(.A(new_n684_), .B(KEYINPUT24), .ZN(new_n685_));
  INV_X1    g0256(.A(new_n685_), .ZN(new_n686_));
  AOI22_X1  g0257(.A1(new_n654_), .A2(G226), .B1(G233), .B2(G335), .ZN(new_n687_));
  INV_X1    g0258(.A(G422), .ZN(new_n688_));
  NAND2_X1  g0259(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g0260(.A1(G233), .A2(G335), .ZN(new_n690_));
  OAI21_X1  g0261(.A(new_n690_), .B1(new_n650_), .B2(new_n608_), .ZN(new_n691_));
  NAND2_X1  g0262(.A1(new_n691_), .A2(G422), .ZN(new_n692_));
  NAND2_X1  g0263(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g0264(.A(new_n693_), .B(KEYINPUT25), .ZN(new_n694_));
  INV_X1    g0265(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g0266(.A1(new_n654_), .A2(G218), .ZN(new_n696_));
  NAND2_X1  g0267(.A1(G225), .A2(G335), .ZN(new_n697_));
  NAND2_X1  g0268(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g0269(.A1(new_n698_), .A2(G468), .ZN(new_n699_));
  NAND3_X1  g0270(.A1(new_n696_), .A2(new_n602_), .A3(new_n697_), .ZN(new_n700_));
  NAND2_X1  g0271(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g0272(.A(new_n701_), .ZN(new_n702_));
  MUX2_X1   g0273(.A(G206), .B(G209), .S(G335), .Z(new_n703_));
  XNOR2_X1  g0274(.A(new_n703_), .B(KEYINPUT26), .ZN(new_n704_));
  XNOR2_X1  g0275(.A(new_n704_), .B(G446), .ZN(new_n705_));
  NOR2_X1   g0276(.A1(new_n630_), .A2(G217), .ZN(new_n706_));
  AOI21_X1  g0277(.A(new_n706_), .B1(new_n617_), .B2(new_n630_), .ZN(new_n707_));
  NOR2_X1   g0278(.A1(new_n707_), .A2(G457), .ZN(new_n708_));
  INV_X1    g0279(.A(new_n708_), .ZN(new_n709_));
  NAND2_X1  g0280(.A1(new_n707_), .A2(G457), .ZN(new_n710_));
  NAND2_X1  g0281(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g0282(.A(new_n711_), .ZN(new_n712_));
  NAND4_X1  g0283(.A1(new_n695_), .A2(new_n702_), .A3(new_n705_), .A4(new_n712_), .ZN(new_n713_));
  NOR2_X1   g0284(.A1(new_n686_), .A2(new_n713_), .ZN(G588));
  MUX2_X1   g0285(.A(G324), .B(G331), .S(G332), .Z(new_n715_));
  XNOR2_X1  g0286(.A(new_n715_), .B(KEYINPUT30), .ZN(new_n716_));
  AND2_X1   g0287(.A1(new_n716_), .A2(G503), .ZN(new_n717_));
  NOR2_X1   g0288(.A1(new_n716_), .A2(G503), .ZN(new_n718_));
  NOR2_X1   g0289(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g0290(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g0291(.A1(G315), .A2(G332), .ZN(new_n721_));
  OR2_X1    g0292(.A1(new_n721_), .A2(KEYINPUT28), .ZN(new_n722_));
  OAI211_X1 g0293(.A(new_n721_), .B(KEYINPUT28), .C1(new_n538_), .C2(G332), .ZN(new_n723_));
  NAND2_X1  g0294(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g0295(.A(new_n724_), .ZN(new_n725_));
  XOR2_X1   g0296(.A(KEYINPUT29), .B(G479), .Z(new_n726_));
  NAND2_X1  g0297(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g0298(.A1(new_n724_), .A2(new_n537_), .ZN(new_n728_));
  NAND2_X1  g0299(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  MUX2_X1   g0300(.A(G316), .B(G323), .S(G332), .Z(new_n730_));
  NOR2_X1   g0301(.A1(new_n730_), .A2(G490), .ZN(new_n731_));
  INV_X1    g0302(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g0303(.A1(new_n730_), .A2(G490), .ZN(new_n733_));
  NAND2_X1  g0304(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g0305(.A1(new_n729_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g0306(.A1(G302), .A2(G332), .ZN(new_n736_));
  INV_X1    g0307(.A(G307), .ZN(new_n737_));
  AOI21_X1  g0308(.A(new_n736_), .B1(new_n737_), .B2(G332), .ZN(new_n738_));
  INV_X1    g0309(.A(new_n738_), .ZN(new_n739_));
  NOR2_X1   g0310(.A1(G293), .A2(G332), .ZN(new_n740_));
  AOI21_X1  g0311(.A(new_n740_), .B1(G593), .B2(G332), .ZN(new_n741_));
  XNOR2_X1  g0312(.A(new_n741_), .B(KEYINPUT27), .ZN(new_n742_));
  NAND3_X1  g0313(.A1(new_n735_), .A2(new_n739_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g0314(.A(G514), .ZN(new_n744_));
  AOI21_X1  g0315(.A(new_n744_), .B1(G611), .B2(G332), .ZN(new_n745_));
  NAND2_X1  g0316(.A1(G611), .A2(G332), .ZN(new_n746_));
  INV_X1    g0317(.A(KEYINPUT31), .ZN(new_n747_));
  XNOR2_X1  g0318(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  AOI21_X1  g0319(.A(new_n745_), .B1(new_n748_), .B2(new_n744_), .ZN(new_n749_));
  INV_X1    g0320(.A(G332), .ZN(new_n750_));
  NAND2_X1  g0321(.A1(new_n750_), .A2(new_n510_), .ZN(new_n751_));
  NAND2_X1  g0322(.A1(G599), .A2(G332), .ZN(new_n752_));
  NAND3_X1  g0323(.A1(new_n751_), .A2(new_n752_), .A3(G523), .ZN(new_n753_));
  INV_X1    g0324(.A(new_n753_), .ZN(new_n754_));
  AOI21_X1  g0325(.A(G523), .B1(new_n751_), .B2(new_n752_), .ZN(new_n755_));
  NOR2_X1   g0326(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g0327(.A1(new_n749_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g0328(.A1(G332), .A2(G358), .ZN(new_n758_));
  INV_X1    g0329(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g0330(.A1(new_n497_), .A2(KEYINPUT7), .ZN(new_n760_));
  INV_X1    g0331(.A(KEYINPUT7), .ZN(new_n761_));
  NAND2_X1  g0332(.A1(new_n761_), .A2(G351), .ZN(new_n762_));
  NAND2_X1  g0333(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g0334(.A(new_n759_), .B1(new_n763_), .B2(new_n750_), .ZN(new_n764_));
  OAI21_X1  g0335(.A(KEYINPUT32), .B1(new_n764_), .B2(G534), .ZN(new_n765_));
  OAI21_X1  g0336(.A(new_n758_), .B1(new_n497_), .B2(G332), .ZN(new_n766_));
  INV_X1    g0337(.A(new_n766_), .ZN(new_n767_));
  NAND2_X1  g0338(.A1(new_n767_), .A2(G534), .ZN(new_n768_));
  OAI21_X1  g0339(.A(new_n758_), .B1(new_n500_), .B2(G332), .ZN(new_n769_));
  INV_X1    g0340(.A(KEYINPUT32), .ZN(new_n770_));
  NAND3_X1  g0341(.A1(new_n769_), .A2(new_n770_), .A3(new_n502_), .ZN(new_n771_));
  NAND3_X1  g0342(.A1(new_n765_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  NOR2_X1   g0343(.A1(G332), .A2(G361), .ZN(new_n773_));
  AOI21_X1  g0344(.A(new_n773_), .B1(G332), .B2(G600), .ZN(new_n774_));
  INV_X1    g0345(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g0346(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  NOR4_X1   g0347(.A1(new_n720_), .A2(new_n743_), .A3(new_n757_), .A4(new_n776_), .ZN(G615));
  NOR4_X1   g0348(.A1(new_n720_), .A2(new_n743_), .A3(new_n757_), .A4(new_n776_), .ZN(G626));
  INV_X1    g0349(.A(new_n629_), .ZN(new_n779_));
  NAND2_X1  g0350(.A1(new_n657_), .A2(new_n672_), .ZN(new_n780_));
  INV_X1    g0351(.A(new_n780_), .ZN(new_n781_));
  AOI22_X1  g0352(.A1(new_n679_), .A2(G400), .B1(new_n677_), .B2(new_n674_), .ZN(new_n782_));
  NAND2_X1  g0353(.A1(new_n669_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g0354(.A1(new_n783_), .A2(new_n643_), .ZN(new_n784_));
  NAND2_X1  g0355(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g0356(.A1(new_n713_), .A2(new_n779_), .A3(new_n785_), .ZN(G632));
  XNOR2_X1  g0357(.A(G361), .B(G369), .ZN(new_n787_));
  XNOR2_X1  g0358(.A(new_n787_), .B(new_n526_), .ZN(new_n788_));
  XNOR2_X1  g0359(.A(G308), .B(G316), .ZN(new_n789_));
  XNOR2_X1  g0360(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g0361(.A(G341), .B(G351), .ZN(new_n791_));
  XNOR2_X1  g0362(.A(G293), .B(G302), .ZN(new_n792_));
  XNOR2_X1  g0363(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g0364(.A(new_n790_), .B(new_n793_), .ZN(G1002));
  XNOR2_X1  g0365(.A(G281), .B(G289), .ZN(new_n795_));
  XNOR2_X1  g0366(.A(new_n795_), .B(KEYINPUT33), .ZN(new_n796_));
  XNOR2_X1  g0367(.A(new_n796_), .B(new_n555_), .ZN(new_n797_));
  XOR2_X1   g0368(.A(G206), .B(G210), .Z(new_n798_));
  XNOR2_X1  g0369(.A(new_n797_), .B(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g0370(.A(G218), .B(G226), .ZN(new_n800_));
  XNOR2_X1  g0371(.A(new_n800_), .B(KEYINPUT34), .ZN(new_n801_));
  XNOR2_X1  g0372(.A(G234), .B(G257), .ZN(new_n802_));
  XNOR2_X1  g0373(.A(new_n802_), .B(new_n659_), .ZN(new_n803_));
  XNOR2_X1  g0374(.A(new_n801_), .B(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g0375(.A(new_n799_), .B(new_n804_), .ZN(G1004));
  AOI21_X1  g0376(.A(new_n602_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n806_));
  NOR2_X1   g0377(.A1(new_n687_), .A2(new_n688_), .ZN(new_n807_));
  AOI21_X1  g0378(.A(new_n806_), .B1(new_n807_), .B2(new_n700_), .ZN(new_n808_));
  AOI21_X1  g0379(.A(new_n708_), .B1(new_n808_), .B2(new_n710_), .ZN(new_n809_));
  NAND2_X1  g0380(.A1(new_n809_), .A2(new_n705_), .ZN(new_n810_));
  AOI21_X1  g0381(.A(new_n558_), .B1(new_n655_), .B2(new_n646_), .ZN(new_n811_));
  NOR3_X1   g0382(.A1(new_n661_), .A2(new_n663_), .A3(KEYINPUT22), .ZN(new_n812_));
  AOI21_X1  g0383(.A(new_n667_), .B1(new_n666_), .B2(new_n660_), .ZN(new_n813_));
  OAI211_X1 g0384(.A(new_n782_), .B(new_n811_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g0385(.A1(new_n645_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g0386(.A1(new_n647_), .A2(new_n649_), .A3(G273), .ZN(new_n816_));
  AOI21_X1  g0387(.A(new_n577_), .B1(new_n816_), .B2(new_n658_), .ZN(new_n817_));
  NAND4_X1  g0388(.A1(new_n639_), .A2(new_n642_), .A3(new_n782_), .A4(new_n817_), .ZN(new_n818_));
  OAI21_X1  g0389(.A(new_n818_), .B1(new_n643_), .B2(new_n680_), .ZN(new_n819_));
  XOR2_X1   g0390(.A(new_n642_), .B(KEYINPUT35), .Z(new_n820_));
  AOI21_X1  g0391(.A(new_n819_), .B1(KEYINPUT36), .B2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g0392(.A1(new_n779_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g0393(.A1(new_n628_), .A2(new_n592_), .ZN(new_n823_));
  AOI21_X1  g0394(.A(KEYINPUT36), .B1(new_n629_), .B2(new_n820_), .ZN(new_n824_));
  NOR4_X1   g0395(.A1(new_n815_), .A2(new_n822_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  OAI221_X1 g0396(.A(new_n810_), .B1(new_n585_), .B2(new_n704_), .C1(new_n825_), .C2(new_n713_), .ZN(G591));
  NOR2_X1   g0397(.A1(new_n738_), .A2(new_n741_), .ZN(new_n827_));
  NOR2_X1   g0398(.A1(new_n724_), .A2(new_n537_), .ZN(new_n828_));
  INV_X1    g0399(.A(KEYINPUT37), .ZN(new_n829_));
  XNOR2_X1  g0400(.A(new_n733_), .B(new_n829_), .ZN(new_n830_));
  INV_X1    g0401(.A(new_n830_), .ZN(new_n831_));
  INV_X1    g0402(.A(new_n729_), .ZN(new_n832_));
  AOI21_X1  g0403(.A(new_n828_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g0404(.A1(new_n766_), .A2(G534), .ZN(new_n834_));
  INV_X1    g0405(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g0406(.A(new_n835_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n836_));
  AOI21_X1  g0407(.A(new_n755_), .B1(new_n836_), .B2(new_n753_), .ZN(new_n837_));
  NAND2_X1  g0408(.A1(new_n837_), .A2(new_n749_), .ZN(new_n838_));
  INV_X1    g0409(.A(new_n748_), .ZN(new_n839_));
  NAND2_X1  g0410(.A1(new_n839_), .A2(G514), .ZN(new_n840_));
  AOI21_X1  g0411(.A(new_n718_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g0412(.A1(new_n841_), .A2(new_n717_), .ZN(new_n842_));
  XOR2_X1   g0413(.A(new_n842_), .B(KEYINPUT38), .Z(new_n843_));
  OAI211_X1 g0414(.A(new_n827_), .B(new_n833_), .C1(new_n843_), .C2(new_n743_), .ZN(G618));
  OAI221_X1 g0415(.A(new_n810_), .B1(new_n585_), .B2(new_n704_), .C1(new_n825_), .C2(new_n713_), .ZN(G621));
  OAI211_X1 g0416(.A(new_n827_), .B(new_n833_), .C1(new_n843_), .C2(new_n743_), .ZN(G629));
  INV_X1    g0417(.A(G4092), .ZN(new_n847_));
  NOR2_X1   g0418(.A1(new_n847_), .A2(G4091), .ZN(new_n848_));
  NAND2_X1  g0419(.A1(new_n848_), .A2(G131), .ZN(new_n849_));
  NOR2_X1   g0420(.A1(G4091), .A2(G4092), .ZN(new_n850_));
  INV_X1    g0421(.A(new_n850_), .ZN(new_n851_));
  OAI21_X1  g0422(.A(new_n849_), .B1(new_n522_), .B2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g0423(.A(new_n774_), .B(G54), .Z(new_n853_));
  INV_X1    g0424(.A(new_n853_), .ZN(new_n854_));
  INV_X1    g0425(.A(G4091), .ZN(new_n855_));
  NOR2_X1   g0426(.A1(new_n855_), .A2(G4092), .ZN(new_n856_));
  AOI21_X1  g0427(.A(new_n852_), .B1(new_n854_), .B2(new_n856_), .ZN(G822));
  AOI22_X1  g0428(.A1(new_n505_), .A2(new_n850_), .B1(G129), .B2(new_n848_), .ZN(new_n858_));
  INV_X1    g0429(.A(new_n856_), .ZN(new_n859_));
  NOR2_X1   g0430(.A1(new_n774_), .A2(G54), .ZN(new_n860_));
  INV_X1    g0431(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g0432(.A(new_n859_), .B1(new_n772_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g0433(.A(new_n862_), .B1(new_n772_), .B2(new_n861_), .ZN(new_n863_));
  NAND2_X1  g0434(.A1(new_n858_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g0435(.A(new_n864_), .ZN(G838));
  OAI21_X1  g0436(.A(new_n855_), .B1(new_n847_), .B2(G117), .ZN(new_n866_));
  AOI21_X1  g0437(.A(new_n866_), .B1(new_n566_), .B2(new_n847_), .ZN(new_n867_));
  XNOR2_X1  g0438(.A(new_n780_), .B(G4), .ZN(new_n868_));
  AOI21_X1  g0439(.A(new_n867_), .B1(new_n868_), .B2(new_n856_), .ZN(G861));
  NAND3_X1  g0440(.A1(new_n772_), .A2(G54), .A3(new_n775_), .ZN(new_n870_));
  OR3_X1    g0441(.A1(new_n720_), .A2(new_n757_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g0442(.A1(new_n843_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g0443(.A(KEYINPUT39), .ZN(new_n873_));
  XNOR2_X1  g0444(.A(new_n872_), .B(new_n873_), .ZN(new_n874_));
  NOR2_X1   g0445(.A1(new_n828_), .A2(new_n738_), .ZN(new_n875_));
  AOI21_X1  g0446(.A(new_n731_), .B1(new_n537_), .B2(new_n724_), .ZN(new_n876_));
  INV_X1    g0447(.A(new_n876_), .ZN(new_n877_));
  INV_X1    g0448(.A(new_n727_), .ZN(new_n878_));
  OAI21_X1  g0449(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g0450(.A(new_n879_), .B(new_n741_), .ZN(new_n880_));
  NAND2_X1  g0451(.A1(new_n874_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g0452(.A1(new_n831_), .A2(new_n832_), .ZN(new_n882_));
  NAND2_X1  g0453(.A1(new_n882_), .A2(new_n875_), .ZN(new_n883_));
  XNOR2_X1  g0454(.A(new_n883_), .B(KEYINPUT40), .ZN(new_n884_));
  INV_X1    g0455(.A(new_n742_), .ZN(new_n885_));
  XNOR2_X1  g0456(.A(new_n884_), .B(new_n885_), .ZN(new_n886_));
  OAI21_X1  g0457(.A(new_n881_), .B1(new_n874_), .B2(new_n886_), .ZN(new_n887_));
  XOR2_X1   g0458(.A(new_n887_), .B(KEYINPUT41), .Z(new_n888_));
  INV_X1    g0459(.A(new_n888_), .ZN(G623));
  OAI21_X1  g0460(.A(G4087), .B1(G11), .B2(G4088), .ZN(new_n890_));
  INV_X1    g0461(.A(G61), .ZN(new_n891_));
  AOI21_X1  g0462(.A(new_n890_), .B1(new_n891_), .B2(G4088), .ZN(new_n892_));
  INV_X1    g0463(.A(G822), .ZN(new_n893_));
  NOR2_X1   g0464(.A1(G4087), .A2(G4088), .ZN(new_n894_));
  AOI21_X1  g0465(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  XOR2_X1   g0466(.A(G861), .B(KEYINPUT42), .Z(new_n896_));
  INV_X1    g0467(.A(new_n896_), .ZN(new_n897_));
  XOR2_X1   g0468(.A(KEYINPUT43), .B(G4087), .Z(new_n898_));
  INV_X1    g0469(.A(new_n898_), .ZN(new_n899_));
  INV_X1    g0470(.A(G4088), .ZN(new_n900_));
  NOR2_X1   g0471(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g0472(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g0473(.A(new_n895_), .B1(new_n897_), .B2(new_n902_), .ZN(G722));
  AOI21_X1  g0474(.A(new_n755_), .B1(new_n753_), .B2(new_n834_), .ZN(new_n904_));
  AOI22_X1  g0475(.A1(new_n749_), .A2(new_n904_), .B1(G514), .B2(new_n839_), .ZN(new_n905_));
  NAND4_X1  g0476(.A1(new_n749_), .A2(new_n756_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n906_));
  NAND2_X1  g0477(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g0478(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g0479(.A(new_n908_), .B1(new_n757_), .B2(new_n870_), .ZN(new_n909_));
  XNOR2_X1  g0480(.A(new_n909_), .B(new_n719_), .ZN(new_n910_));
  NOR2_X1   g0481(.A1(new_n535_), .A2(G4092), .ZN(new_n911_));
  OAI21_X1  g0482(.A(new_n855_), .B1(new_n847_), .B2(G52), .ZN(new_n912_));
  OAI22_X1  g0483(.A1(new_n910_), .A2(new_n859_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g0484(.A(new_n913_), .B(KEYINPUT44), .ZN(new_n914_));
  INV_X1    g0485(.A(new_n914_), .ZN(G832));
  INV_X1    g0486(.A(new_n772_), .ZN(new_n916_));
  NOR3_X1   g0487(.A1(new_n916_), .A2(new_n755_), .A3(new_n860_), .ZN(new_n917_));
  NOR2_X1   g0488(.A1(new_n917_), .A2(new_n904_), .ZN(new_n918_));
  XNOR2_X1  g0489(.A(new_n918_), .B(new_n749_), .ZN(new_n919_));
  NAND2_X1  g0490(.A1(new_n524_), .A2(new_n847_), .ZN(new_n920_));
  INV_X1    g0491(.A(G130), .ZN(new_n921_));
  AOI21_X1  g0492(.A(G4091), .B1(new_n921_), .B2(G4092), .ZN(new_n922_));
  AOI22_X1  g0493(.A1(new_n919_), .A2(new_n856_), .B1(new_n920_), .B2(new_n922_), .ZN(G834));
  XNOR2_X1  g0494(.A(new_n766_), .B(G534), .ZN(new_n924_));
  OAI211_X1 g0495(.A(new_n870_), .B(new_n834_), .C1(new_n775_), .C2(new_n924_), .ZN(new_n925_));
  XOR2_X1   g0496(.A(new_n756_), .B(KEYINPUT45), .Z(new_n926_));
  XNOR2_X1  g0497(.A(new_n925_), .B(new_n926_), .ZN(new_n927_));
  NOR2_X1   g0498(.A1(new_n927_), .A2(new_n859_), .ZN(new_n928_));
  OAI21_X1  g0499(.A(new_n855_), .B1(new_n847_), .B2(G119), .ZN(new_n929_));
  AOI21_X1  g0500(.A(new_n929_), .B1(new_n512_), .B2(new_n847_), .ZN(new_n930_));
  NOR2_X1   g0501(.A1(new_n928_), .A2(new_n930_), .ZN(G836));
  OAI21_X1  g0502(.A(G4090), .B1(G11), .B2(G4089), .ZN(new_n932_));
  AOI21_X1  g0503(.A(new_n932_), .B1(new_n891_), .B2(G4089), .ZN(new_n933_));
  NOR2_X1   g0504(.A1(G4089), .A2(G4090), .ZN(new_n934_));
  AOI21_X1  g0505(.A(new_n933_), .B1(new_n893_), .B2(new_n934_), .ZN(new_n935_));
  XOR2_X1   g0506(.A(KEYINPUT46), .B(G4090), .Z(new_n936_));
  INV_X1    g0507(.A(new_n936_), .ZN(new_n937_));
  INV_X1    g0508(.A(G4089), .ZN(new_n938_));
  NOR2_X1   g0509(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  INV_X1    g0510(.A(new_n939_), .ZN(new_n940_));
  OAI21_X1  g0511(.A(new_n935_), .B1(new_n897_), .B2(new_n940_), .ZN(G859));
  INV_X1    g0512(.A(G4), .ZN(new_n942_));
  NOR2_X1   g0513(.A1(new_n780_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g0514(.A1(new_n943_), .A2(new_n784_), .ZN(new_n944_));
  OAI21_X1  g0515(.A(KEYINPUT48), .B1(new_n814_), .B2(new_n643_), .ZN(new_n945_));
  AND2_X1   g0516(.A1(new_n639_), .A2(new_n642_), .ZN(new_n946_));
  NAND2_X1  g0517(.A1(new_n674_), .A2(new_n677_), .ZN(new_n947_));
  NAND2_X1  g0518(.A1(new_n680_), .A2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g0519(.A(new_n948_), .B1(new_n664_), .B2(new_n668_), .ZN(new_n949_));
  INV_X1    g0520(.A(KEYINPUT48), .ZN(new_n950_));
  NAND4_X1  g0521(.A1(new_n946_), .A2(new_n949_), .A3(new_n950_), .A4(new_n811_), .ZN(new_n951_));
  INV_X1    g0522(.A(new_n817_), .ZN(new_n952_));
  NOR2_X1   g0523(.A1(new_n952_), .A2(new_n948_), .ZN(new_n953_));
  INV_X1    g0524(.A(KEYINPUT47), .ZN(new_n954_));
  NAND3_X1  g0525(.A1(new_n946_), .A2(new_n953_), .A3(new_n954_), .ZN(new_n955_));
  NAND2_X1  g0526(.A1(new_n818_), .A2(KEYINPUT47), .ZN(new_n956_));
  AOI22_X1  g0527(.A1(new_n945_), .A2(new_n951_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g0528(.A1(new_n944_), .A2(new_n957_), .ZN(new_n958_));
  OR2_X1    g0529(.A1(new_n958_), .A2(KEYINPUT49), .ZN(new_n959_));
  NOR2_X1   g0530(.A1(new_n643_), .A2(new_n680_), .ZN(new_n960_));
  NOR2_X1   g0531(.A1(new_n820_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g0532(.A1(new_n958_), .A2(KEYINPUT49), .ZN(new_n962_));
  NAND3_X1  g0533(.A1(new_n959_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  XNOR2_X1  g0534(.A(new_n963_), .B(new_n779_), .ZN(new_n964_));
  AND2_X1   g0535(.A1(new_n964_), .A2(new_n856_), .ZN(new_n965_));
  OAI21_X1  g0536(.A(new_n855_), .B1(new_n847_), .B2(G122), .ZN(new_n966_));
  AOI21_X1  g0537(.A(new_n966_), .B1(new_n600_), .B2(new_n847_), .ZN(new_n967_));
  NOR2_X1   g0538(.A1(new_n965_), .A2(new_n967_), .ZN(G871));
  NAND2_X1  g0539(.A1(new_n943_), .A2(new_n949_), .ZN(new_n969_));
  INV_X1    g0540(.A(KEYINPUT50), .ZN(new_n970_));
  NAND4_X1  g0541(.A1(new_n669_), .A2(new_n970_), .A3(new_n782_), .A4(new_n811_), .ZN(new_n971_));
  AOI21_X1  g0542(.A(new_n681_), .B1(new_n817_), .B2(new_n675_), .ZN(new_n972_));
  NAND2_X1  g0543(.A1(new_n814_), .A2(KEYINPUT50), .ZN(new_n973_));
  NAND4_X1  g0544(.A1(new_n969_), .A2(new_n971_), .A3(new_n972_), .A4(new_n973_), .ZN(new_n974_));
  XNOR2_X1  g0545(.A(new_n974_), .B(new_n946_), .ZN(new_n975_));
  OR2_X1    g0546(.A1(new_n975_), .A2(new_n859_), .ZN(new_n976_));
  NAND3_X1  g0547(.A1(new_n570_), .A2(new_n847_), .A3(new_n573_), .ZN(new_n977_));
  INV_X1    g0548(.A(KEYINPUT51), .ZN(new_n978_));
  AOI22_X1  g0549(.A1(new_n977_), .A2(new_n978_), .B1(G128), .B2(G4092), .ZN(new_n979_));
  OAI21_X1  g0550(.A(new_n979_), .B1(new_n978_), .B2(new_n977_), .ZN(new_n980_));
  NAND2_X1  g0551(.A1(new_n980_), .A2(new_n855_), .ZN(new_n981_));
  NAND2_X1  g0552(.A1(new_n976_), .A2(new_n981_), .ZN(new_n982_));
  INV_X1    g0553(.A(new_n982_), .ZN(G873));
  AOI22_X1  g0554(.A1(new_n654_), .A2(G273), .B1(G280), .B2(G335), .ZN(new_n984_));
  OAI21_X1  g0555(.A(new_n660_), .B1(new_n984_), .B2(G411), .ZN(new_n985_));
  NAND2_X1  g0556(.A1(new_n985_), .A2(new_n811_), .ZN(new_n986_));
  OR2_X1    g0557(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n987_));
  NAND2_X1  g0558(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n988_));
  NAND3_X1  g0559(.A1(new_n986_), .A2(new_n987_), .A3(new_n988_), .ZN(new_n989_));
  AOI21_X1  g0560(.A(new_n989_), .B1(new_n943_), .B2(new_n669_), .ZN(new_n990_));
  XNOR2_X1  g0561(.A(new_n782_), .B(KEYINPUT53), .ZN(new_n991_));
  XNOR2_X1  g0562(.A(new_n990_), .B(new_n991_), .ZN(new_n992_));
  NOR2_X1   g0563(.A1(new_n992_), .A2(new_n859_), .ZN(new_n993_));
  OAI21_X1  g0564(.A(new_n855_), .B1(new_n847_), .B2(G127), .ZN(new_n994_));
  AOI21_X1  g0565(.A(new_n994_), .B1(new_n557_), .B2(new_n847_), .ZN(new_n995_));
  NOR2_X1   g0566(.A1(new_n993_), .A2(new_n995_), .ZN(G875));
  NOR2_X1   g0567(.A1(new_n943_), .A2(new_n811_), .ZN(new_n997_));
  XNOR2_X1  g0568(.A(new_n997_), .B(new_n669_), .ZN(new_n998_));
  AND2_X1   g0569(.A1(new_n998_), .A2(new_n856_), .ZN(new_n999_));
  NOR2_X1   g0570(.A1(new_n580_), .A2(G4092), .ZN(new_n1000_));
  INV_X1    g0571(.A(new_n1000_), .ZN(new_n1001_));
  OR2_X1    g0572(.A1(new_n1001_), .A2(KEYINPUT54), .ZN(new_n1002_));
  AOI22_X1  g0573(.A1(new_n1001_), .A2(KEYINPUT54), .B1(G126), .B2(G4092), .ZN(new_n1003_));
  AOI21_X1  g0574(.A(G4091), .B1(new_n1002_), .B2(new_n1003_), .ZN(new_n1004_));
  NOR2_X1   g0575(.A1(new_n999_), .A2(new_n1004_), .ZN(G877));
  XNOR2_X1  g0576(.A(new_n748_), .B(KEYINPUT56), .ZN(new_n1006_));
  XNOR2_X1  g0577(.A(new_n1006_), .B(new_n775_), .ZN(new_n1007_));
  XNOR2_X1  g0578(.A(new_n738_), .B(new_n741_), .ZN(new_n1008_));
  XNOR2_X1  g0579(.A(new_n1007_), .B(new_n1008_), .ZN(new_n1009_));
  NAND2_X1  g0580(.A1(new_n751_), .A2(new_n752_), .ZN(new_n1010_));
  XNOR2_X1  g0581(.A(new_n716_), .B(new_n1010_), .ZN(new_n1011_));
  XNOR2_X1  g0582(.A(new_n1011_), .B(new_n769_), .ZN(new_n1012_));
  MUX2_X1   g0583(.A(G369), .B(G372), .S(G332), .Z(new_n1013_));
  XNOR2_X1  g0584(.A(new_n1013_), .B(KEYINPUT55), .ZN(new_n1014_));
  XNOR2_X1  g0585(.A(new_n1012_), .B(new_n1014_), .ZN(new_n1015_));
  XNOR2_X1  g0586(.A(new_n1009_), .B(new_n1015_), .ZN(new_n1016_));
  XNOR2_X1  g0587(.A(new_n1016_), .B(new_n730_), .ZN(new_n1017_));
  XNOR2_X1  g0588(.A(new_n1017_), .B(new_n724_), .ZN(G998));
  XNOR2_X1  g0589(.A(new_n691_), .B(KEYINPUT57), .ZN(new_n1019_));
  XNOR2_X1  g0590(.A(new_n1019_), .B(new_n704_), .ZN(new_n1020_));
  MUX2_X1   g0591(.A(G289), .B(G292), .S(G335), .Z(new_n1021_));
  XNOR2_X1  g0592(.A(new_n1020_), .B(new_n1021_), .ZN(new_n1022_));
  XOR2_X1   g0593(.A(new_n628_), .B(new_n707_), .Z(new_n1023_));
  XNOR2_X1  g0594(.A(new_n1022_), .B(new_n1023_), .ZN(new_n1024_));
  NAND2_X1  g0595(.A1(new_n670_), .A2(new_n671_), .ZN(new_n1025_));
  XOR2_X1   g0596(.A(new_n679_), .B(new_n665_), .Z(new_n1026_));
  XNOR2_X1  g0597(.A(new_n1025_), .B(new_n1026_), .ZN(new_n1027_));
  XNOR2_X1  g0598(.A(new_n1024_), .B(new_n1027_), .ZN(new_n1028_));
  XNOR2_X1  g0599(.A(new_n698_), .B(KEYINPUT58), .ZN(new_n1029_));
  NOR2_X1   g0600(.A1(new_n633_), .A2(new_n638_), .ZN(new_n1030_));
  XNOR2_X1  g0601(.A(new_n1029_), .B(new_n1030_), .ZN(new_n1031_));
  XNOR2_X1  g0602(.A(new_n1028_), .B(new_n1031_), .ZN(G1000));
  NOR2_X1   g0603(.A1(new_n785_), .A2(new_n779_), .ZN(new_n1033_));
  AOI21_X1  g0604(.A(new_n942_), .B1(new_n1033_), .B2(KEYINPUT59), .ZN(new_n1034_));
  OAI21_X1  g0605(.A(new_n1034_), .B1(KEYINPUT59), .B2(new_n1033_), .ZN(new_n1035_));
  NAND2_X1  g0606(.A1(new_n1035_), .A2(new_n825_), .ZN(new_n1036_));
  XNOR2_X1  g0607(.A(new_n1036_), .B(KEYINPUT60), .ZN(new_n1037_));
  XNOR2_X1  g0608(.A(new_n1037_), .B(new_n695_), .ZN(new_n1038_));
  XNOR2_X1  g0609(.A(new_n1037_), .B(KEYINPUT61), .ZN(new_n1039_));
  XNOR2_X1  g0610(.A(new_n809_), .B(new_n705_), .ZN(new_n1040_));
  AND2_X1   g0611(.A1(new_n689_), .A2(new_n700_), .ZN(new_n1041_));
  NOR2_X1   g0612(.A1(new_n1041_), .A2(new_n806_), .ZN(new_n1042_));
  NAND2_X1  g0613(.A1(new_n1042_), .A2(new_n710_), .ZN(new_n1043_));
  NAND2_X1  g0614(.A1(new_n1043_), .A2(new_n709_), .ZN(new_n1044_));
  INV_X1    g0615(.A(new_n705_), .ZN(new_n1045_));
  XNOR2_X1  g0616(.A(new_n1044_), .B(new_n1045_), .ZN(new_n1046_));
  OAI22_X1  g0617(.A1(new_n1039_), .A2(new_n1040_), .B1(new_n1037_), .B2(new_n1046_), .ZN(new_n1047_));
  XNOR2_X1  g0618(.A(new_n711_), .B(new_n808_), .ZN(new_n1048_));
  XNOR2_X1  g0619(.A(new_n1042_), .B(new_n711_), .ZN(new_n1049_));
  OAI22_X1  g0620(.A1(new_n1039_), .A2(new_n1048_), .B1(new_n1037_), .B2(new_n1049_), .ZN(new_n1050_));
  AOI211_X1 g0621(.A(new_n1038_), .B(new_n1047_), .C1(KEYINPUT62), .C2(new_n1050_), .ZN(new_n1051_));
  AOI21_X1  g0622(.A(new_n807_), .B1(new_n1039_), .B2(new_n689_), .ZN(new_n1052_));
  XNOR2_X1  g0623(.A(new_n1052_), .B(new_n701_), .ZN(new_n1053_));
  OAI211_X1 g0624(.A(new_n1051_), .B(new_n1053_), .C1(KEYINPUT62), .C2(new_n1050_), .ZN(new_n1054_));
  XNOR2_X1  g0625(.A(new_n1054_), .B(KEYINPUT63), .ZN(new_n1055_));
  NOR2_X1   g0626(.A1(new_n998_), .A2(new_n868_), .ZN(new_n1056_));
  NAND3_X1  g0627(.A1(new_n975_), .A2(new_n1056_), .A3(new_n992_), .ZN(new_n1057_));
  NOR3_X1   g0628(.A1(new_n1055_), .A2(new_n964_), .A3(new_n1057_), .ZN(G575));
  NAND2_X1  g0629(.A1(new_n874_), .A2(new_n731_), .ZN(new_n1059_));
  OAI21_X1  g0630(.A(new_n1059_), .B1(new_n831_), .B2(new_n874_), .ZN(new_n1060_));
  XNOR2_X1  g0631(.A(new_n1060_), .B(new_n729_), .ZN(new_n1061_));
  NAND2_X1  g0632(.A1(new_n874_), .A2(new_n735_), .ZN(new_n1062_));
  NAND2_X1  g0633(.A1(new_n1062_), .A2(new_n833_), .ZN(new_n1063_));
  XNOR2_X1  g0634(.A(new_n1063_), .B(new_n739_), .ZN(new_n1064_));
  XOR2_X1   g0635(.A(new_n874_), .B(new_n734_), .Z(new_n1065_));
  NAND4_X1  g0636(.A1(G623), .A2(new_n1061_), .A3(new_n1064_), .A4(new_n1065_), .ZN(new_n1066_));
  XOR2_X1   g0637(.A(new_n1066_), .B(KEYINPUT64), .Z(new_n1067_));
  NOR3_X1   g0638(.A1(new_n919_), .A2(new_n916_), .A3(new_n854_), .ZN(new_n1068_));
  AND4_X1   g0639(.A1(new_n910_), .A2(new_n1067_), .A3(new_n927_), .A4(new_n1068_), .ZN(G585));
  INV_X1    g0640(.A(G137), .ZN(new_n1070_));
  INV_X1    g0641(.A(G1689), .ZN(new_n1071_));
  NOR2_X1   g0642(.A1(new_n1071_), .A2(G1690), .ZN(new_n1072_));
  NAND2_X1  g0643(.A1(new_n896_), .A2(new_n1072_), .ZN(new_n1073_));
  XOR2_X1   g0644(.A(new_n1073_), .B(KEYINPUT65), .Z(new_n1074_));
  OAI21_X1  g0645(.A(G1690), .B1(G182), .B2(G1689), .ZN(new_n1075_));
  INV_X1    g0646(.A(G185), .ZN(new_n1076_));
  AOI21_X1  g0647(.A(new_n1075_), .B1(new_n1076_), .B2(G1689), .ZN(new_n1077_));
  NOR2_X1   g0648(.A1(G1689), .A2(G1690), .ZN(new_n1078_));
  AOI21_X1  g0649(.A(new_n1077_), .B1(new_n893_), .B2(new_n1078_), .ZN(new_n1079_));
  AOI21_X1  g0650(.A(new_n1070_), .B1(new_n1074_), .B2(new_n1079_), .ZN(G661));
  INV_X1    g0651(.A(G1691), .ZN(new_n1081_));
  NOR2_X1   g0652(.A1(new_n1081_), .A2(G1694), .ZN(new_n1082_));
  INV_X1    g0653(.A(new_n1082_), .ZN(new_n1083_));
  NOR2_X1   g0654(.A1(new_n897_), .A2(new_n1083_), .ZN(new_n1084_));
  NOR2_X1   g0655(.A1(G822), .A2(G1694), .ZN(new_n1085_));
  NAND2_X1  g0656(.A1(new_n1085_), .A2(KEYINPUT66), .ZN(new_n1086_));
  INV_X1    g0657(.A(new_n1086_), .ZN(new_n1087_));
  OAI21_X1  g0658(.A(G1694), .B1(G182), .B2(G1691), .ZN(new_n1088_));
  OAI21_X1  g0659(.A(new_n1088_), .B1(new_n1085_), .B2(KEYINPUT66), .ZN(new_n1089_));
  OAI21_X1  g0660(.A(new_n1081_), .B1(new_n1087_), .B2(new_n1089_), .ZN(new_n1090_));
  OAI21_X1  g0661(.A(new_n1090_), .B1(new_n1076_), .B2(new_n1088_), .ZN(new_n1091_));
  OAI21_X1  g0662(.A(G137), .B1(new_n1084_), .B2(new_n1091_), .ZN(new_n1092_));
  XOR2_X1   g0663(.A(new_n1092_), .B(KEYINPUT67), .Z(G693));
  OR2_X1    g0664(.A1(G43), .A2(G4088), .ZN(new_n1094_));
  OAI211_X1 g0665(.A(new_n1094_), .B(G4087), .C1(G37), .C2(new_n900_), .ZN(new_n1095_));
  NOR2_X1   g0666(.A1(new_n899_), .A2(G4088), .ZN(new_n1096_));
  INV_X1    g0667(.A(new_n1096_), .ZN(new_n1097_));
  OAI221_X1 g0668(.A(new_n1095_), .B1(G871), .B2(new_n902_), .C1(G832), .C2(new_n1097_), .ZN(G747));
  INV_X1    g0669(.A(G834), .ZN(new_n1099_));
  NAND2_X1  g0670(.A1(new_n1099_), .A2(new_n1096_), .ZN(new_n1100_));
  NOR2_X1   g0671(.A1(new_n900_), .A2(G20), .ZN(new_n1101_));
  OAI21_X1  g0672(.A(G4087), .B1(G76), .B2(G4088), .ZN(new_n1102_));
  OAI221_X1 g0673(.A(new_n1100_), .B1(new_n1101_), .B2(new_n1102_), .C1(G873), .C2(new_n902_), .ZN(G752));
  INV_X1    g0674(.A(G17), .ZN(new_n1104_));
  NAND2_X1  g0675(.A1(new_n1104_), .A2(G4088), .ZN(new_n1105_));
  OAI211_X1 g0676(.A(new_n1105_), .B(G4087), .C1(G73), .C2(G4088), .ZN(new_n1106_));
  OAI221_X1 g0677(.A(new_n1106_), .B1(G836), .B2(new_n1097_), .C1(G875), .C2(new_n902_), .ZN(G757));
  NAND2_X1  g0678(.A1(new_n864_), .A2(new_n894_), .ZN(new_n1108_));
  NOR2_X1   g0679(.A1(new_n900_), .A2(G70), .ZN(new_n1109_));
  OAI21_X1  g0680(.A(G4087), .B1(G67), .B2(G4088), .ZN(new_n1110_));
  OAI221_X1 g0681(.A(new_n1108_), .B1(new_n1109_), .B2(new_n1110_), .C1(G877), .C2(new_n902_), .ZN(G762));
  NOR2_X1   g0682(.A1(new_n937_), .A2(G4089), .ZN(new_n1112_));
  NAND2_X1  g0683(.A1(new_n914_), .A2(new_n1112_), .ZN(new_n1113_));
  XNOR2_X1  g0684(.A(new_n1113_), .B(KEYINPUT68), .ZN(new_n1114_));
  NOR2_X1   g0685(.A1(new_n938_), .A2(G37), .ZN(new_n1115_));
  OAI21_X1  g0686(.A(G4090), .B1(G43), .B2(G4089), .ZN(new_n1116_));
  OAI221_X1 g0687(.A(new_n1114_), .B1(new_n940_), .B2(G871), .C1(new_n1115_), .C2(new_n1116_), .ZN(G787));
  NAND2_X1  g0688(.A1(new_n1099_), .A2(new_n1112_), .ZN(new_n1118_));
  NOR2_X1   g0689(.A1(new_n938_), .A2(G20), .ZN(new_n1119_));
  OAI21_X1  g0690(.A(G4090), .B1(G76), .B2(G4089), .ZN(new_n1120_));
  OAI221_X1 g0691(.A(new_n1118_), .B1(new_n1119_), .B2(new_n1120_), .C1(G873), .C2(new_n940_), .ZN(G792));
  NAND2_X1  g0692(.A1(new_n1104_), .A2(G4089), .ZN(new_n1122_));
  OAI211_X1 g0693(.A(new_n1122_), .B(G4090), .C1(G73), .C2(G4089), .ZN(new_n1123_));
  INV_X1    g0694(.A(new_n1112_), .ZN(new_n1124_));
  OAI221_X1 g0695(.A(new_n1123_), .B1(G836), .B2(new_n1124_), .C1(G875), .C2(new_n940_), .ZN(G797));
  NAND2_X1  g0696(.A1(new_n864_), .A2(new_n934_), .ZN(new_n1126_));
  NOR2_X1   g0697(.A1(new_n938_), .A2(G70), .ZN(new_n1127_));
  OAI21_X1  g0698(.A(G4090), .B1(G67), .B2(G4089), .ZN(new_n1128_));
  OAI221_X1 g0699(.A(new_n1126_), .B1(new_n1127_), .B2(new_n1128_), .C1(G877), .C2(new_n940_), .ZN(new_n1129_));
  XNOR2_X1  g0700(.A(new_n1129_), .B(KEYINPUT69), .ZN(G802));
  INV_X1    g0701(.A(G871), .ZN(new_n1131_));
  NAND2_X1  g0702(.A1(new_n1131_), .A2(new_n1072_), .ZN(new_n1132_));
  NAND3_X1  g0703(.A1(G170), .A2(G1689), .A3(G1690), .ZN(new_n1133_));
  INV_X1    g0704(.A(G200), .ZN(new_n1134_));
  INV_X1    g0705(.A(G1690), .ZN(new_n1135_));
  OAI21_X1  g0706(.A(KEYINPUT70), .B1(new_n1134_), .B2(new_n1135_), .ZN(new_n1136_));
  NAND2_X1  g0707(.A1(new_n1136_), .A2(new_n1071_), .ZN(new_n1137_));
  NOR3_X1   g0708(.A1(new_n1134_), .A2(new_n1135_), .A3(KEYINPUT70), .ZN(new_n1138_));
  OAI21_X1  g0709(.A(new_n1133_), .B1(new_n1137_), .B2(new_n1138_), .ZN(new_n1139_));
  AOI21_X1  g0710(.A(new_n1139_), .B1(new_n914_), .B2(new_n1078_), .ZN(new_n1140_));
  AOI21_X1  g0711(.A(new_n1070_), .B1(new_n1132_), .B2(new_n1140_), .ZN(G642));
  OAI21_X1  g0712(.A(new_n1072_), .B1(new_n999_), .B2(new_n1004_), .ZN(new_n1142_));
  OAI21_X1  g0713(.A(G1690), .B1(G188), .B2(G1689), .ZN(new_n1143_));
  INV_X1    g0714(.A(G158), .ZN(new_n1144_));
  AOI21_X1  g0715(.A(new_n1143_), .B1(new_n1144_), .B2(G1689), .ZN(new_n1145_));
  AOI21_X1  g0716(.A(new_n1145_), .B1(new_n864_), .B2(new_n1078_), .ZN(new_n1146_));
  AOI21_X1  g0717(.A(new_n1070_), .B1(new_n1142_), .B2(new_n1146_), .ZN(G664));
  INV_X1    g0718(.A(G875), .ZN(new_n1148_));
  NAND2_X1  g0719(.A1(new_n1148_), .A2(new_n1072_), .ZN(new_n1149_));
  OAI21_X1  g0720(.A(G1690), .B1(G155), .B2(G1689), .ZN(new_n1150_));
  INV_X1    g0721(.A(G152), .ZN(new_n1151_));
  AOI21_X1  g0722(.A(new_n1150_), .B1(new_n1151_), .B2(G1689), .ZN(new_n1152_));
  INV_X1    g0723(.A(G836), .ZN(new_n1153_));
  AOI21_X1  g0724(.A(new_n1152_), .B1(new_n1153_), .B2(new_n1078_), .ZN(new_n1154_));
  AOI21_X1  g0725(.A(new_n1070_), .B1(new_n1149_), .B2(new_n1154_), .ZN(G667));
  NAND2_X1  g0726(.A1(new_n982_), .A2(new_n1072_), .ZN(new_n1156_));
  XOR2_X1   g0727(.A(new_n1156_), .B(KEYINPUT71), .Z(new_n1157_));
  OAI21_X1  g0728(.A(G1690), .B1(G149), .B2(G1689), .ZN(new_n1158_));
  INV_X1    g0729(.A(G146), .ZN(new_n1159_));
  AOI21_X1  g0730(.A(new_n1158_), .B1(new_n1159_), .B2(G1689), .ZN(new_n1160_));
  AOI21_X1  g0731(.A(new_n1160_), .B1(new_n1099_), .B2(new_n1078_), .ZN(new_n1161_));
  AOI21_X1  g0732(.A(new_n1070_), .B1(new_n1157_), .B2(new_n1161_), .ZN(G670));
  NAND2_X1  g0733(.A1(new_n1131_), .A2(new_n1082_), .ZN(new_n1163_));
  OAI21_X1  g0734(.A(G1694), .B1(G200), .B2(G1691), .ZN(new_n1164_));
  INV_X1    g0735(.A(G170), .ZN(new_n1165_));
  AOI21_X1  g0736(.A(new_n1164_), .B1(new_n1165_), .B2(G1691), .ZN(new_n1166_));
  NOR2_X1   g0737(.A1(G1691), .A2(G1694), .ZN(new_n1167_));
  AOI21_X1  g0738(.A(new_n1166_), .B1(new_n914_), .B2(new_n1167_), .ZN(new_n1168_));
  AOI21_X1  g0739(.A(new_n1070_), .B1(new_n1163_), .B2(new_n1168_), .ZN(G676));
  NOR2_X1   g0740(.A1(G877), .A2(new_n1083_), .ZN(new_n1170_));
  XNOR2_X1  g0741(.A(new_n1170_), .B(KEYINPUT72), .ZN(new_n1171_));
  OAI21_X1  g0742(.A(G1694), .B1(G188), .B2(G1691), .ZN(new_n1172_));
  AOI21_X1  g0743(.A(new_n1172_), .B1(new_n1144_), .B2(G1691), .ZN(new_n1173_));
  AOI21_X1  g0744(.A(new_n1173_), .B1(new_n864_), .B2(new_n1167_), .ZN(new_n1174_));
  AOI21_X1  g0745(.A(new_n1070_), .B1(new_n1171_), .B2(new_n1174_), .ZN(G696));
  NAND2_X1  g0746(.A1(new_n1148_), .A2(new_n1082_), .ZN(new_n1176_));
  OAI21_X1  g0747(.A(G1694), .B1(G155), .B2(G1691), .ZN(new_n1177_));
  AOI21_X1  g0748(.A(new_n1177_), .B1(new_n1151_), .B2(G1691), .ZN(new_n1178_));
  AOI21_X1  g0749(.A(new_n1178_), .B1(new_n1153_), .B2(new_n1167_), .ZN(new_n1179_));
  AOI21_X1  g0750(.A(new_n1070_), .B1(new_n1176_), .B2(new_n1179_), .ZN(G699));
  NAND2_X1  g0751(.A1(new_n982_), .A2(new_n1082_), .ZN(new_n1181_));
  OAI21_X1  g0752(.A(G1694), .B1(G149), .B2(G1691), .ZN(new_n1182_));
  AOI21_X1  g0753(.A(new_n1182_), .B1(new_n1159_), .B2(G1691), .ZN(new_n1183_));
  AOI21_X1  g0754(.A(new_n1183_), .B1(new_n1099_), .B2(new_n1167_), .ZN(new_n1184_));
  AOI21_X1  g0755(.A(new_n1070_), .B1(new_n1181_), .B2(new_n1184_), .ZN(G702));
  NAND2_X1  g0756(.A1(G135), .A2(G4115), .ZN(new_n1186_));
  NOR2_X1   g0757(.A1(new_n516_), .A2(G3717), .ZN(new_n1187_));
  INV_X1    g0758(.A(G3724), .ZN(new_n1188_));
  INV_X1    g0759(.A(G123), .ZN(new_n1189_));
  INV_X1    g0760(.A(G3717), .ZN(new_n1190_));
  OAI21_X1  g0761(.A(new_n1188_), .B1(new_n1189_), .B2(new_n1190_), .ZN(new_n1191_));
  OAI21_X1  g0762(.A(new_n1186_), .B1(new_n1187_), .B2(new_n1191_), .ZN(new_n1192_));
  NAND2_X1  g0763(.A1(new_n888_), .A2(G3717), .ZN(new_n1193_));
  XNOR2_X1  g0764(.A(new_n741_), .B(G132), .ZN(new_n1194_));
  AOI21_X1  g0765(.A(new_n1188_), .B1(new_n1194_), .B2(new_n1190_), .ZN(new_n1195_));
  AOI21_X1  g0766(.A(new_n1192_), .B1(new_n1193_), .B2(new_n1195_), .ZN(G818));
  XOR2_X1   g0767(.A(new_n888_), .B(new_n1194_), .Z(G813));
  OAI21_X1  g0768(.A(new_n855_), .B1(new_n847_), .B2(G123), .ZN(new_n1198_));
  AOI21_X1  g0769(.A(new_n1198_), .B1(new_n516_), .B2(new_n847_), .ZN(new_n1199_));
  AOI21_X1  g0770(.A(new_n1199_), .B1(new_n888_), .B2(new_n856_), .ZN(G824));
  NOR2_X1   g0771(.A1(new_n1064_), .A2(new_n859_), .ZN(new_n1201_));
  OAI21_X1  g0772(.A(new_n855_), .B1(new_n847_), .B2(G121), .ZN(new_n1202_));
  AOI21_X1  g0773(.A(new_n1202_), .B1(new_n519_), .B2(new_n847_), .ZN(new_n1203_));
  NOR2_X1   g0774(.A1(new_n1201_), .A2(new_n1203_), .ZN(G826));
  NOR2_X1   g0775(.A1(new_n1061_), .A2(new_n859_), .ZN(new_n1205_));
  OAI21_X1  g0776(.A(new_n855_), .B1(new_n847_), .B2(G116), .ZN(new_n1206_));
  AOI21_X1  g0777(.A(new_n1206_), .B1(new_n543_), .B2(new_n847_), .ZN(new_n1207_));
  NOR2_X1   g0778(.A1(new_n1205_), .A2(new_n1207_), .ZN(G828));
  NAND2_X1  g0779(.A1(new_n549_), .A2(new_n546_), .ZN(new_n1209_));
  NOR2_X1   g0780(.A1(new_n1209_), .A2(G4092), .ZN(new_n1210_));
  OAI21_X1  g0781(.A(new_n855_), .B1(new_n847_), .B2(G112), .ZN(new_n1211_));
  OAI22_X1  g0782(.A1(new_n1065_), .A2(new_n859_), .B1(new_n1210_), .B2(new_n1211_), .ZN(new_n1212_));
  XOR2_X1   g0783(.A(new_n1212_), .B(KEYINPUT73), .Z(new_n1213_));
  INV_X1    g0784(.A(new_n1213_), .ZN(G830));
  NAND3_X1  g0785(.A1(G601), .A2(G245), .A3(G559), .ZN(new_n1215_));
  OR3_X1    g0786(.A1(G1002), .A2(G847), .A3(new_n1215_), .ZN(new_n1216_));
  NOR4_X1   g0787(.A1(G998), .A2(G1004), .A3(G1000), .A4(new_n1216_), .ZN(G854));
  AND2_X1   g0788(.A1(new_n1047_), .A2(new_n856_), .ZN(new_n1218_));
  OAI21_X1  g0789(.A(new_n855_), .B1(new_n847_), .B2(G115), .ZN(new_n1219_));
  AOI21_X1  g0790(.A(new_n1219_), .B1(new_n591_), .B2(new_n847_), .ZN(new_n1220_));
  NOR2_X1   g0791(.A1(new_n1218_), .A2(new_n1220_), .ZN(G863));
  AND2_X1   g0792(.A1(new_n1050_), .A2(new_n856_), .ZN(new_n1222_));
  OAI21_X1  g0793(.A(new_n855_), .B1(new_n847_), .B2(G114), .ZN(new_n1223_));
  AOI21_X1  g0794(.A(new_n1223_), .B1(new_n625_), .B2(new_n847_), .ZN(new_n1224_));
  NOR2_X1   g0795(.A1(new_n1222_), .A2(new_n1224_), .ZN(G865));
  OR3_X1    g0796(.A1(new_n1053_), .A2(KEYINPUT74), .A3(new_n859_), .ZN(new_n1226_));
  NAND2_X1  g0797(.A1(new_n607_), .A2(new_n847_), .ZN(new_n1227_));
  OAI211_X1 g0798(.A(new_n1227_), .B(new_n855_), .C1(G53), .C2(new_n847_), .ZN(new_n1228_));
  OAI21_X1  g0799(.A(KEYINPUT74), .B1(new_n1053_), .B2(new_n859_), .ZN(new_n1229_));
  NAND3_X1  g0800(.A1(new_n1226_), .A2(new_n1228_), .A3(new_n1229_), .ZN(new_n1230_));
  INV_X1    g0801(.A(new_n1230_), .ZN(G867));
  NAND2_X1  g0802(.A1(new_n613_), .A2(new_n847_), .ZN(new_n1232_));
  OAI211_X1 g0803(.A(new_n1232_), .B(new_n855_), .C1(G113), .C2(new_n847_), .ZN(new_n1233_));
  INV_X1    g0804(.A(new_n1038_), .ZN(new_n1234_));
  OAI21_X1  g0805(.A(new_n1233_), .B1(new_n1234_), .B2(new_n859_), .ZN(new_n1235_));
  XNOR2_X1  g0806(.A(new_n1235_), .B(KEYINPUT75), .ZN(new_n1236_));
  INV_X1    g0807(.A(new_n1236_), .ZN(G869));
  NAND3_X1  g0808(.A1(new_n938_), .A2(G109), .A3(G4090), .ZN(new_n1238_));
  XNOR2_X1  g0809(.A(new_n1238_), .B(KEYINPUT76), .ZN(new_n1239_));
  AND3_X1   g0810(.A1(G106), .A2(G4089), .A3(G4090), .ZN(new_n1240_));
  INV_X1    g0811(.A(G863), .ZN(new_n1241_));
  AOI211_X1 g0812(.A(new_n1239_), .B(new_n1240_), .C1(new_n1241_), .C2(new_n939_), .ZN(new_n1242_));
  OAI21_X1  g0813(.A(new_n1242_), .B1(G824), .B2(new_n1124_), .ZN(G712));
  OR2_X1    g0814(.A1(G109), .A2(G4088), .ZN(new_n1244_));
  OAI211_X1 g0815(.A(new_n1244_), .B(G4087), .C1(G106), .C2(new_n900_), .ZN(new_n1245_));
  OAI221_X1 g0816(.A(new_n1245_), .B1(new_n902_), .B2(G863), .C1(G824), .C2(new_n1097_), .ZN(G727));
  OAI21_X1  g0817(.A(G4087), .B1(G46), .B2(G4088), .ZN(new_n1247_));
  INV_X1    g0818(.A(G49), .ZN(new_n1248_));
  AOI21_X1  g0819(.A(new_n1247_), .B1(new_n1248_), .B2(G4088), .ZN(new_n1249_));
  INV_X1    g0820(.A(G865), .ZN(new_n1250_));
  AOI21_X1  g0821(.A(new_n1249_), .B1(new_n1250_), .B2(new_n901_), .ZN(new_n1251_));
  OAI21_X1  g0822(.A(new_n1251_), .B1(G826), .B2(new_n1097_), .ZN(G732));
  OAI21_X1  g0823(.A(G4087), .B1(G100), .B2(G4088), .ZN(new_n1253_));
  INV_X1    g0824(.A(G103), .ZN(new_n1254_));
  AOI21_X1  g0825(.A(new_n1253_), .B1(new_n1254_), .B2(G4088), .ZN(new_n1255_));
  AOI21_X1  g0826(.A(new_n1255_), .B1(new_n1230_), .B2(new_n901_), .ZN(new_n1256_));
  OAI21_X1  g0827(.A(new_n1256_), .B1(new_n1097_), .B2(G828), .ZN(G737));
  OAI21_X1  g0828(.A(G4087), .B1(G91), .B2(G4088), .ZN(new_n1258_));
  INV_X1    g0829(.A(G40), .ZN(new_n1259_));
  AOI21_X1  g0830(.A(new_n1258_), .B1(new_n1259_), .B2(G4088), .ZN(new_n1260_));
  AOI21_X1  g0831(.A(new_n1260_), .B1(new_n1236_), .B2(new_n901_), .ZN(new_n1261_));
  OAI21_X1  g0832(.A(new_n1261_), .B1(G830), .B2(new_n1097_), .ZN(G742));
  OAI21_X1  g0833(.A(G4090), .B1(G46), .B2(G4089), .ZN(new_n1263_));
  AOI21_X1  g0834(.A(new_n1263_), .B1(new_n1248_), .B2(G4089), .ZN(new_n1264_));
  AOI21_X1  g0835(.A(new_n1264_), .B1(new_n1250_), .B2(new_n939_), .ZN(new_n1265_));
  OAI21_X1  g0836(.A(new_n1265_), .B1(G826), .B2(new_n1124_), .ZN(G772));
  OAI21_X1  g0837(.A(G4090), .B1(G100), .B2(G4089), .ZN(new_n1267_));
  AOI21_X1  g0838(.A(new_n1267_), .B1(new_n1254_), .B2(G4089), .ZN(new_n1268_));
  AOI21_X1  g0839(.A(new_n1268_), .B1(new_n1230_), .B2(new_n939_), .ZN(new_n1269_));
  OAI21_X1  g0840(.A(new_n1269_), .B1(new_n1124_), .B2(G828), .ZN(G777));
  OAI21_X1  g0841(.A(G4090), .B1(G91), .B2(G4089), .ZN(new_n1271_));
  AOI21_X1  g0842(.A(new_n1271_), .B1(new_n1259_), .B2(G4089), .ZN(new_n1272_));
  AOI21_X1  g0843(.A(new_n1272_), .B1(new_n1236_), .B2(new_n939_), .ZN(new_n1273_));
  OAI21_X1  g0844(.A(new_n1273_), .B1(G830), .B2(new_n1124_), .ZN(G782));
  NAND2_X1  g0845(.A1(new_n1213_), .A2(new_n1078_), .ZN(new_n1275_));
  OAI21_X1  g0846(.A(G1690), .B1(G203), .B2(G1689), .ZN(new_n1276_));
  INV_X1    g0847(.A(G173), .ZN(new_n1277_));
  AOI21_X1  g0848(.A(new_n1276_), .B1(new_n1277_), .B2(G1689), .ZN(new_n1278_));
  AOI21_X1  g0849(.A(new_n1278_), .B1(new_n1236_), .B2(new_n1072_), .ZN(new_n1279_));
  AOI21_X1  g0850(.A(new_n1070_), .B1(new_n1275_), .B2(new_n1279_), .ZN(G645));
  OAI21_X1  g0851(.A(G1690), .B1(G197), .B2(G1689), .ZN(new_n1281_));
  INV_X1    g0852(.A(G167), .ZN(new_n1282_));
  AOI21_X1  g0853(.A(new_n1281_), .B1(new_n1282_), .B2(G1689), .ZN(new_n1283_));
  AOI21_X1  g0854(.A(new_n1283_), .B1(new_n1230_), .B2(new_n1072_), .ZN(new_n1284_));
  OAI21_X1  g0855(.A(new_n1078_), .B1(new_n1205_), .B2(new_n1207_), .ZN(new_n1285_));
  AOI21_X1  g0856(.A(new_n1070_), .B1(new_n1284_), .B2(new_n1285_), .ZN(G648));
  OAI21_X1  g0857(.A(new_n1078_), .B1(new_n1201_), .B2(new_n1203_), .ZN(new_n1287_));
  OAI21_X1  g0858(.A(G1690), .B1(G194), .B2(G1689), .ZN(new_n1288_));
  INV_X1    g0859(.A(G164), .ZN(new_n1289_));
  AOI21_X1  g0860(.A(new_n1288_), .B1(new_n1289_), .B2(G1689), .ZN(new_n1290_));
  AOI21_X1  g0861(.A(new_n1290_), .B1(new_n1250_), .B2(new_n1072_), .ZN(new_n1291_));
  AOI21_X1  g0862(.A(new_n1070_), .B1(new_n1287_), .B2(new_n1291_), .ZN(G651));
  OR3_X1    g0863(.A1(G824), .A2(G1689), .A3(G1690), .ZN(new_n1293_));
  OAI21_X1  g0864(.A(G1690), .B1(G191), .B2(G1689), .ZN(new_n1294_));
  INV_X1    g0865(.A(G161), .ZN(new_n1295_));
  AOI21_X1  g0866(.A(new_n1294_), .B1(new_n1295_), .B2(G1689), .ZN(new_n1296_));
  AOI21_X1  g0867(.A(new_n1296_), .B1(new_n1241_), .B2(new_n1072_), .ZN(new_n1297_));
  AOI21_X1  g0868(.A(new_n1070_), .B1(new_n1293_), .B2(new_n1297_), .ZN(G654));
  NAND2_X1  g0869(.A1(new_n1213_), .A2(new_n1167_), .ZN(new_n1299_));
  OAI21_X1  g0870(.A(G1694), .B1(G203), .B2(G1691), .ZN(new_n1300_));
  AOI21_X1  g0871(.A(new_n1300_), .B1(new_n1277_), .B2(G1691), .ZN(new_n1301_));
  XNOR2_X1  g0872(.A(new_n1301_), .B(KEYINPUT77), .ZN(new_n1302_));
  AOI21_X1  g0873(.A(new_n1302_), .B1(new_n1236_), .B2(new_n1082_), .ZN(new_n1303_));
  AOI21_X1  g0874(.A(new_n1070_), .B1(new_n1299_), .B2(new_n1303_), .ZN(G679));
  NAND2_X1  g0875(.A1(new_n1282_), .A2(G1691), .ZN(new_n1305_));
  OAI211_X1 g0876(.A(new_n1305_), .B(G1694), .C1(G197), .C2(G1691), .ZN(new_n1306_));
  OAI21_X1  g0877(.A(new_n1306_), .B1(G867), .B2(new_n1083_), .ZN(new_n1307_));
  INV_X1    g0878(.A(new_n1167_), .ZN(new_n1308_));
  NOR2_X1   g0879(.A1(G828), .A2(new_n1308_), .ZN(new_n1309_));
  OAI21_X1  g0880(.A(G137), .B1(new_n1307_), .B2(new_n1309_), .ZN(new_n1310_));
  XNOR2_X1  g0881(.A(new_n1310_), .B(KEYINPUT78), .ZN(G682));
  NAND2_X1  g0882(.A1(new_n1289_), .A2(G1691), .ZN(new_n1312_));
  OAI211_X1 g0883(.A(new_n1312_), .B(G1694), .C1(G194), .C2(G1691), .ZN(new_n1313_));
  OAI21_X1  g0884(.A(new_n1313_), .B1(G826), .B2(new_n1308_), .ZN(new_n1314_));
  INV_X1    g0885(.A(KEYINPUT79), .ZN(new_n1315_));
  OAI22_X1  g0886(.A1(new_n1314_), .A2(new_n1315_), .B1(new_n1083_), .B2(G865), .ZN(new_n1316_));
  AND2_X1   g0887(.A1(new_n1314_), .A2(new_n1315_), .ZN(new_n1317_));
  OAI21_X1  g0888(.A(G137), .B1(new_n1316_), .B2(new_n1317_), .ZN(new_n1318_));
  NAND2_X1  g0889(.A1(new_n1318_), .A2(KEYINPUT80), .ZN(new_n1319_));
  INV_X1    g0890(.A(KEYINPUT80), .ZN(new_n1320_));
  OAI211_X1 g0891(.A(new_n1320_), .B(G137), .C1(new_n1316_), .C2(new_n1317_), .ZN(new_n1321_));
  NAND2_X1  g0892(.A1(new_n1319_), .A2(new_n1321_), .ZN(G685));
  NOR2_X1   g0893(.A1(G824), .A2(G1694), .ZN(new_n1323_));
  AOI21_X1  g0894(.A(G1691), .B1(new_n1323_), .B2(KEYINPUT81), .ZN(new_n1324_));
  OAI21_X1  g0895(.A(new_n1324_), .B1(KEYINPUT81), .B2(new_n1323_), .ZN(new_n1325_));
  NAND2_X1  g0896(.A1(new_n1295_), .A2(G1691), .ZN(new_n1326_));
  OAI211_X1 g0897(.A(new_n1326_), .B(G1694), .C1(G191), .C2(G1691), .ZN(new_n1327_));
  NOR2_X1   g0898(.A1(G863), .A2(new_n1083_), .ZN(new_n1328_));
  OAI21_X1  g0899(.A(new_n1327_), .B1(new_n1328_), .B2(KEYINPUT82), .ZN(new_n1329_));
  AOI21_X1  g0900(.A(new_n1329_), .B1(KEYINPUT82), .B2(new_n1328_), .ZN(new_n1330_));
  AOI21_X1  g0901(.A(new_n1070_), .B1(new_n1325_), .B2(new_n1330_), .ZN(G688));
  OAI21_X1  g0902(.A(G4092), .B1(G120), .B2(G4091), .ZN(new_n1332_));
  XOR2_X1   g0903(.A(new_n1332_), .B(KEYINPUT98), .Z(new_n1333_));
  NAND3_X1  g0904(.A1(G248), .A2(G324), .A3(G503), .ZN(new_n1334_));
  XNOR2_X1  g0905(.A(new_n1334_), .B(KEYINPUT95), .ZN(new_n1335_));
  NAND3_X1  g0906(.A1(new_n526_), .A2(G251), .A3(G503), .ZN(new_n1336_));
  AOI21_X1  g0907(.A(G503), .B1(new_n526_), .B2(G254), .ZN(new_n1337_));
  OAI21_X1  g0908(.A(new_n1337_), .B1(new_n514_), .B2(new_n526_), .ZN(new_n1338_));
  NAND3_X1  g0909(.A1(new_n1335_), .A2(new_n1336_), .A3(new_n1338_), .ZN(new_n1339_));
  XNOR2_X1  g0910(.A(new_n1339_), .B(KEYINPUT96), .ZN(new_n1340_));
  MUX2_X1   g0911(.A(new_n514_), .B(G248), .S(G514), .Z(new_n1341_));
  XNOR2_X1  g0912(.A(new_n1340_), .B(new_n1341_), .ZN(new_n1342_));
  OR2_X1    g0913(.A1(new_n1342_), .A2(new_n522_), .ZN(new_n1343_));
  NAND3_X1  g0914(.A1(new_n510_), .A2(G251), .A3(G523), .ZN(new_n1344_));
  XNOR2_X1  g0915(.A(new_n1344_), .B(KEYINPUT93), .ZN(new_n1345_));
  NAND3_X1  g0916(.A1(G248), .A2(G341), .A3(G523), .ZN(new_n1346_));
  NOR2_X1   g0917(.A1(new_n514_), .A2(new_n510_), .ZN(new_n1347_));
  INV_X1    g0918(.A(G523), .ZN(new_n1348_));
  OAI21_X1  g0919(.A(new_n1348_), .B1(new_n540_), .B2(G341), .ZN(new_n1349_));
  OAI211_X1 g0920(.A(new_n1345_), .B(new_n1346_), .C1(new_n1347_), .C2(new_n1349_), .ZN(new_n1350_));
  XNOR2_X1  g0921(.A(new_n1350_), .B(KEYINPUT94), .ZN(new_n1351_));
  AOI21_X1  g0922(.A(G534), .B1(new_n497_), .B2(G254), .ZN(new_n1352_));
  OAI21_X1  g0923(.A(new_n1352_), .B1(new_n514_), .B2(new_n497_), .ZN(new_n1353_));
  AOI22_X1  g0924(.A1(new_n500_), .A2(G251), .B1(G248), .B2(G351), .ZN(new_n1354_));
  OAI21_X1  g0925(.A(new_n1353_), .B1(new_n1354_), .B2(new_n502_), .ZN(new_n1355_));
  XNOR2_X1  g0926(.A(new_n1351_), .B(new_n1355_), .ZN(new_n1356_));
  NOR2_X1   g0927(.A1(new_n1343_), .A2(new_n1356_), .ZN(new_n1357_));
  XNOR2_X1  g0928(.A(new_n1357_), .B(KEYINPUT97), .ZN(new_n1358_));
  NAND2_X1  g0929(.A1(new_n1342_), .A2(new_n522_), .ZN(new_n1359_));
  NAND3_X1  g0930(.A1(new_n1343_), .A2(new_n1356_), .A3(new_n1359_), .ZN(new_n1360_));
  OAI211_X1 g0931(.A(new_n1358_), .B(new_n1360_), .C1(new_n1356_), .C2(new_n1359_), .ZN(new_n1361_));
  XNOR2_X1  g0932(.A(new_n1209_), .B(new_n543_), .ZN(new_n1362_));
  XOR2_X1   g0933(.A(new_n519_), .B(new_n515_), .Z(new_n1363_));
  XNOR2_X1  g0934(.A(new_n1362_), .B(new_n1363_), .ZN(new_n1364_));
  XNOR2_X1  g0935(.A(new_n1361_), .B(new_n1364_), .ZN(new_n1365_));
  AOI21_X1  g0936(.A(new_n1333_), .B1(new_n1365_), .B2(new_n850_), .ZN(new_n1366_));
  INV_X1    g0937(.A(new_n749_), .ZN(new_n1367_));
  NAND3_X1  g0938(.A1(new_n749_), .A2(new_n756_), .A3(new_n772_), .ZN(new_n1368_));
  AND2_X1   g0939(.A1(new_n905_), .A2(new_n1368_), .ZN(new_n1369_));
  NAND3_X1  g0940(.A1(new_n765_), .A2(new_n502_), .A3(new_n771_), .ZN(new_n1370_));
  NOR3_X1   g0941(.A1(new_n1370_), .A2(KEYINPUT88), .A3(new_n904_), .ZN(new_n1371_));
  INV_X1    g0942(.A(new_n755_), .ZN(new_n1372_));
  AOI21_X1  g0943(.A(new_n1371_), .B1(new_n1372_), .B2(new_n1370_), .ZN(new_n1373_));
  XNOR2_X1  g0944(.A(new_n1369_), .B(new_n1373_), .ZN(new_n1374_));
  XNOR2_X1  g0945(.A(new_n772_), .B(new_n774_), .ZN(new_n1375_));
  XNOR2_X1  g0946(.A(new_n1374_), .B(new_n1375_), .ZN(new_n1376_));
  OR2_X1    g0947(.A1(new_n1376_), .A2(new_n719_), .ZN(new_n1377_));
  NAND2_X1  g0948(.A1(new_n1376_), .A2(new_n719_), .ZN(new_n1378_));
  AOI21_X1  g0949(.A(new_n1367_), .B1(new_n1377_), .B2(new_n1378_), .ZN(new_n1379_));
  INV_X1    g0950(.A(new_n1379_), .ZN(new_n1380_));
  INV_X1    g0951(.A(KEYINPUT89), .ZN(new_n1381_));
  NAND2_X1  g0952(.A1(new_n1377_), .A2(new_n1381_), .ZN(new_n1382_));
  NAND3_X1  g0953(.A1(new_n1377_), .A2(new_n1367_), .A3(new_n1378_), .ZN(new_n1383_));
  NAND4_X1  g0954(.A1(new_n1380_), .A2(new_n756_), .A3(new_n1382_), .A4(new_n1383_), .ZN(new_n1384_));
  NAND2_X1  g0955(.A1(new_n1382_), .A2(new_n756_), .ZN(new_n1385_));
  INV_X1    g0956(.A(new_n1383_), .ZN(new_n1386_));
  OAI21_X1  g0957(.A(new_n1385_), .B1(new_n1386_), .B2(new_n1379_), .ZN(new_n1387_));
  NAND3_X1  g0958(.A1(new_n1384_), .A2(new_n1387_), .A3(G2174), .ZN(new_n1388_));
  OR3_X1    g0959(.A1(new_n904_), .A2(KEYINPUT83), .A3(new_n774_), .ZN(new_n1389_));
  OAI21_X1  g0960(.A(KEYINPUT83), .B1(new_n904_), .B2(new_n774_), .ZN(new_n1390_));
  NAND3_X1  g0961(.A1(new_n767_), .A2(new_n753_), .A3(new_n502_), .ZN(new_n1391_));
  NOR2_X1   g0962(.A1(new_n775_), .A2(new_n755_), .ZN(new_n1392_));
  AOI22_X1  g0963(.A1(new_n1389_), .A2(new_n1390_), .B1(new_n1391_), .B2(new_n1392_), .ZN(new_n1393_));
  NAND2_X1  g0964(.A1(new_n1393_), .A2(new_n836_), .ZN(new_n1394_));
  INV_X1    g0965(.A(new_n1394_), .ZN(new_n1395_));
  NOR2_X1   g0966(.A1(new_n1393_), .A2(new_n836_), .ZN(new_n1396_));
  OAI21_X1  g0967(.A(new_n907_), .B1(new_n1395_), .B2(new_n1396_), .ZN(new_n1397_));
  INV_X1    g0968(.A(KEYINPUT84), .ZN(new_n1398_));
  NAND2_X1  g0969(.A1(new_n1397_), .A2(new_n1398_), .ZN(new_n1399_));
  XNOR2_X1  g0970(.A(new_n1393_), .B(new_n836_), .ZN(new_n1400_));
  NAND3_X1  g0971(.A1(new_n1400_), .A2(KEYINPUT84), .A3(new_n907_), .ZN(new_n1401_));
  NAND2_X1  g0972(.A1(new_n1399_), .A2(new_n1401_), .ZN(new_n1402_));
  NOR2_X1   g0973(.A1(new_n904_), .A2(new_n774_), .ZN(new_n1403_));
  AOI21_X1  g0974(.A(new_n1403_), .B1(new_n837_), .B2(new_n774_), .ZN(new_n1404_));
  OAI211_X1 g0975(.A(new_n908_), .B(new_n1394_), .C1(new_n1404_), .C2(new_n836_), .ZN(new_n1405_));
  INV_X1    g0976(.A(new_n1405_), .ZN(new_n1406_));
  OAI21_X1  g0977(.A(new_n774_), .B1(new_n1402_), .B2(new_n1406_), .ZN(new_n1407_));
  NAND4_X1  g0978(.A1(new_n1405_), .A2(new_n1399_), .A3(new_n775_), .A4(new_n1401_), .ZN(new_n1408_));
  NAND3_X1  g0979(.A1(new_n1407_), .A2(KEYINPUT85), .A3(new_n1408_), .ZN(new_n1409_));
  INV_X1    g0980(.A(KEYINPUT85), .ZN(new_n1410_));
  OAI211_X1 g0981(.A(new_n1410_), .B(new_n774_), .C1(new_n1402_), .C2(new_n1406_), .ZN(new_n1411_));
  NAND3_X1  g0982(.A1(new_n1409_), .A2(new_n916_), .A3(new_n1411_), .ZN(new_n1412_));
  OAI21_X1  g0983(.A(new_n1394_), .B1(new_n1404_), .B2(new_n836_), .ZN(new_n1413_));
  NOR2_X1   g0984(.A1(new_n1413_), .A2(new_n908_), .ZN(new_n1414_));
  NAND2_X1  g0985(.A1(new_n1400_), .A2(new_n1369_), .ZN(new_n1415_));
  NAND2_X1  g0986(.A1(new_n1415_), .A2(new_n774_), .ZN(new_n1416_));
  OR3_X1    g0987(.A1(new_n1414_), .A2(KEYINPUT86), .A3(new_n1416_), .ZN(new_n1417_));
  OAI21_X1  g0988(.A(KEYINPUT86), .B1(new_n1414_), .B2(new_n1416_), .ZN(new_n1418_));
  NAND4_X1  g0989(.A1(new_n1417_), .A2(new_n772_), .A3(new_n1408_), .A4(new_n1418_), .ZN(new_n1419_));
  AOI21_X1  g0990(.A(new_n719_), .B1(new_n1412_), .B2(new_n1419_), .ZN(new_n1420_));
  INV_X1    g0991(.A(new_n1420_), .ZN(new_n1421_));
  INV_X1    g0992(.A(KEYINPUT87), .ZN(new_n1422_));
  NAND3_X1  g0993(.A1(new_n1412_), .A2(new_n719_), .A3(new_n1419_), .ZN(new_n1423_));
  NAND4_X1  g0994(.A1(new_n1421_), .A2(new_n1422_), .A3(new_n756_), .A4(new_n1423_), .ZN(new_n1424_));
  NAND2_X1  g0995(.A1(new_n1424_), .A2(new_n1367_), .ZN(new_n1425_));
  NAND3_X1  g0996(.A1(new_n1409_), .A2(new_n772_), .A3(new_n1411_), .ZN(new_n1426_));
  NAND4_X1  g0997(.A1(new_n1417_), .A2(new_n916_), .A3(new_n1408_), .A4(new_n1418_), .ZN(new_n1427_));
  NAND3_X1  g0998(.A1(new_n1426_), .A2(new_n720_), .A3(new_n1427_), .ZN(new_n1428_));
  NAND2_X1  g0999(.A1(new_n1423_), .A2(new_n1428_), .ZN(new_n1429_));
  INV_X1    g1000(.A(new_n756_), .ZN(new_n1430_));
  NAND2_X1  g1001(.A1(new_n1429_), .A2(new_n1430_), .ZN(new_n1431_));
  INV_X1    g1002(.A(new_n1423_), .ZN(new_n1432_));
  NOR2_X1   g1003(.A1(new_n1432_), .A2(new_n1420_), .ZN(new_n1433_));
  AOI21_X1  g1004(.A(new_n1422_), .B1(new_n1433_), .B2(new_n756_), .ZN(new_n1434_));
  AOI21_X1  g1005(.A(new_n1425_), .B1(new_n1431_), .B2(new_n1434_), .ZN(new_n1435_));
  NAND3_X1  g1006(.A1(new_n1423_), .A2(new_n1428_), .A3(new_n756_), .ZN(new_n1436_));
  OAI211_X1 g1007(.A(new_n749_), .B(new_n1436_), .C1(new_n1433_), .C2(new_n756_), .ZN(new_n1437_));
  INV_X1    g1008(.A(G2174), .ZN(new_n1438_));
  NAND2_X1  g1009(.A1(new_n1437_), .A2(new_n1438_), .ZN(new_n1439_));
  OAI21_X1  g1010(.A(new_n1388_), .B1(new_n1435_), .B2(new_n1439_), .ZN(new_n1440_));
  OR4_X1    g1011(.A1(new_n1438_), .A2(new_n720_), .A3(new_n757_), .A4(new_n776_), .ZN(new_n1441_));
  AND2_X1   g1012(.A1(new_n843_), .A2(new_n1441_), .ZN(new_n1442_));
  XNOR2_X1  g1013(.A(new_n879_), .B(new_n734_), .ZN(new_n1443_));
  NAND2_X1  g1014(.A1(new_n727_), .A2(new_n731_), .ZN(new_n1444_));
  AOI21_X1  g1015(.A(new_n832_), .B1(new_n877_), .B2(new_n1444_), .ZN(new_n1445_));
  XNOR2_X1  g1016(.A(new_n1443_), .B(new_n1445_), .ZN(new_n1446_));
  NAND2_X1  g1017(.A1(new_n1446_), .A2(new_n885_), .ZN(new_n1447_));
  OAI21_X1  g1018(.A(new_n1447_), .B1(new_n741_), .B2(new_n1446_), .ZN(new_n1448_));
  NOR2_X1   g1019(.A1(new_n1442_), .A2(new_n1448_), .ZN(new_n1449_));
  INV_X1    g1020(.A(new_n828_), .ZN(new_n1450_));
  AOI21_X1  g1021(.A(new_n830_), .B1(new_n729_), .B2(new_n1450_), .ZN(new_n1451_));
  INV_X1    g1022(.A(KEYINPUT90), .ZN(new_n1452_));
  NAND2_X1  g1023(.A1(new_n1451_), .A2(new_n1452_), .ZN(new_n1453_));
  OAI21_X1  g1024(.A(KEYINPUT90), .B1(new_n831_), .B2(new_n878_), .ZN(new_n1454_));
  OAI21_X1  g1025(.A(new_n1453_), .B1(new_n1451_), .B2(new_n1454_), .ZN(new_n1455_));
  NAND2_X1  g1026(.A1(new_n1455_), .A2(new_n832_), .ZN(new_n1456_));
  OAI211_X1 g1027(.A(new_n1453_), .B(new_n729_), .C1(new_n1451_), .C2(new_n1454_), .ZN(new_n1457_));
  AOI21_X1  g1028(.A(new_n734_), .B1(new_n1456_), .B2(new_n1457_), .ZN(new_n1458_));
  INV_X1    g1029(.A(new_n1458_), .ZN(new_n1459_));
  NAND3_X1  g1030(.A1(new_n1456_), .A2(new_n734_), .A3(new_n1457_), .ZN(new_n1460_));
  NAND4_X1  g1031(.A1(new_n1459_), .A2(new_n882_), .A3(new_n875_), .A4(new_n1460_), .ZN(new_n1461_));
  INV_X1    g1032(.A(new_n1460_), .ZN(new_n1462_));
  OAI21_X1  g1033(.A(new_n883_), .B1(new_n1462_), .B2(new_n1458_), .ZN(new_n1463_));
  NAND3_X1  g1034(.A1(new_n1461_), .A2(new_n1463_), .A3(new_n741_), .ZN(new_n1464_));
  INV_X1    g1035(.A(KEYINPUT91), .ZN(new_n1465_));
  OR2_X1    g1036(.A1(new_n1464_), .A2(new_n1465_), .ZN(new_n1466_));
  NAND2_X1  g1037(.A1(new_n1461_), .A2(new_n1463_), .ZN(new_n1467_));
  NAND2_X1  g1038(.A1(new_n1467_), .A2(new_n742_), .ZN(new_n1468_));
  INV_X1    g1039(.A(KEYINPUT92), .ZN(new_n1469_));
  NAND2_X1  g1040(.A1(new_n1468_), .A2(new_n1469_), .ZN(new_n1470_));
  NAND2_X1  g1041(.A1(new_n1464_), .A2(new_n1465_), .ZN(new_n1471_));
  NAND3_X1  g1042(.A1(new_n1467_), .A2(KEYINPUT92), .A3(new_n742_), .ZN(new_n1472_));
  NAND4_X1  g1043(.A1(new_n1466_), .A2(new_n1470_), .A3(new_n1471_), .A4(new_n1472_), .ZN(new_n1473_));
  AOI21_X1  g1044(.A(new_n1449_), .B1(new_n1473_), .B2(new_n1442_), .ZN(new_n1474_));
  NOR2_X1   g1045(.A1(new_n1474_), .A2(new_n739_), .ZN(new_n1475_));
  AOI211_X1 g1046(.A(new_n738_), .B(new_n1449_), .C1(new_n1473_), .C2(new_n1442_), .ZN(new_n1476_));
  NOR2_X1   g1047(.A1(new_n1475_), .A2(new_n1476_), .ZN(new_n1477_));
  NAND2_X1  g1048(.A1(new_n1440_), .A2(new_n1477_), .ZN(new_n1478_));
  NAND3_X1  g1049(.A1(new_n1421_), .A2(new_n756_), .A3(new_n1423_), .ZN(new_n1479_));
  AND3_X1   g1050(.A1(new_n1479_), .A2(new_n1431_), .A3(KEYINPUT87), .ZN(new_n1480_));
  OAI211_X1 g1051(.A(new_n1438_), .B(new_n1437_), .C1(new_n1480_), .C2(new_n1425_), .ZN(new_n1481_));
  INV_X1    g1052(.A(new_n1477_), .ZN(new_n1482_));
  NAND3_X1  g1053(.A1(new_n1481_), .A2(new_n1388_), .A3(new_n1482_), .ZN(new_n1483_));
  NAND2_X1  g1054(.A1(new_n1478_), .A2(new_n1483_), .ZN(new_n1484_));
  INV_X1    g1055(.A(new_n1484_), .ZN(new_n1485_));
  OAI21_X1  g1056(.A(new_n1366_), .B1(new_n1485_), .B2(new_n859_), .ZN(G843));
  OAI21_X1  g1057(.A(G4092), .B1(G118), .B2(G4091), .ZN(new_n1487_));
  NOR2_X1   g1058(.A1(new_n604_), .A2(new_n518_), .ZN(new_n1488_));
  XNOR2_X1  g1059(.A(new_n1488_), .B(KEYINPUT119), .ZN(new_n1489_));
  AOI21_X1  g1060(.A(G468), .B1(G218), .B2(G242), .ZN(new_n1490_));
  INV_X1    g1061(.A(new_n1490_), .ZN(new_n1491_));
  OAI22_X1  g1062(.A1(new_n1491_), .A2(KEYINPUT118), .B1(G218), .B2(new_n540_), .ZN(new_n1492_));
  AND2_X1   g1063(.A1(new_n1491_), .A2(KEYINPUT118), .ZN(new_n1493_));
  OAI221_X1 g1064(.A(new_n1489_), .B1(new_n1492_), .B2(new_n1493_), .C1(new_n545_), .C2(new_n606_), .ZN(new_n1494_));
  XNOR2_X1  g1065(.A(new_n590_), .B(new_n1494_), .ZN(new_n1495_));
  AOI21_X1  g1066(.A(G422), .B1(new_n608_), .B2(G254), .ZN(new_n1496_));
  OAI21_X1  g1067(.A(new_n1496_), .B1(new_n608_), .B2(new_n514_), .ZN(new_n1497_));
  OAI221_X1 g1068(.A(new_n1497_), .B1(new_n518_), .B2(new_n612_), .C1(new_n545_), .C2(new_n611_), .ZN(new_n1498_));
  XNOR2_X1  g1069(.A(new_n1495_), .B(new_n1498_), .ZN(new_n1499_));
  OAI21_X1  g1070(.A(new_n577_), .B1(new_n514_), .B2(new_n659_), .ZN(new_n1500_));
  OR2_X1    g1071(.A1(new_n1500_), .A2(KEYINPUT115), .ZN(new_n1501_));
  NAND2_X1  g1072(.A1(new_n1500_), .A2(KEYINPUT115), .ZN(new_n1502_));
  OAI211_X1 g1073(.A(new_n1501_), .B(new_n1502_), .C1(new_n540_), .C2(G273), .ZN(new_n1503_));
  NAND3_X1  g1074(.A1(new_n659_), .A2(G251), .A3(G411), .ZN(new_n1504_));
  NAND3_X1  g1075(.A1(G248), .A2(G273), .A3(G411), .ZN(new_n1505_));
  AND2_X1   g1076(.A1(new_n1505_), .A2(KEYINPUT116), .ZN(new_n1506_));
  NOR2_X1   g1077(.A1(new_n1505_), .A2(KEYINPUT116), .ZN(new_n1507_));
  OAI211_X1 g1078(.A(new_n1503_), .B(new_n1504_), .C1(new_n1506_), .C2(new_n1507_), .ZN(new_n1508_));
  NAND3_X1  g1079(.A1(G248), .A2(G281), .A3(G374), .ZN(new_n1509_));
  XNOR2_X1  g1080(.A(new_n1509_), .B(KEYINPUT117), .ZN(new_n1510_));
  NAND3_X1  g1081(.A1(new_n559_), .A2(G251), .A3(G374), .ZN(new_n1511_));
  AOI21_X1  g1082(.A(G374), .B1(new_n559_), .B2(G254), .ZN(new_n1512_));
  OAI21_X1  g1083(.A(new_n1512_), .B1(new_n514_), .B2(new_n559_), .ZN(new_n1513_));
  NAND3_X1  g1084(.A1(new_n1510_), .A2(new_n1511_), .A3(new_n1513_), .ZN(new_n1514_));
  XNOR2_X1  g1085(.A(new_n1508_), .B(new_n1514_), .ZN(new_n1515_));
  NAND2_X1  g1086(.A1(G234), .A2(G242), .ZN(new_n1516_));
  OAI211_X1 g1087(.A(new_n1516_), .B(new_n592_), .C1(G234), .C2(new_n540_), .ZN(new_n1517_));
  OAI221_X1 g1088(.A(new_n1517_), .B1(new_n518_), .B2(new_n595_), .C1(new_n593_), .C2(new_n545_), .ZN(new_n1518_));
  XOR2_X1   g1089(.A(new_n1515_), .B(new_n1518_), .Z(new_n1519_));
  XNOR2_X1  g1090(.A(new_n1499_), .B(new_n1519_), .ZN(new_n1520_));
  NAND3_X1  g1091(.A1(new_n568_), .A2(G251), .A3(G389), .ZN(new_n1521_));
  XOR2_X1   g1092(.A(new_n1521_), .B(KEYINPUT114), .Z(new_n1522_));
  NAND3_X1  g1093(.A1(G248), .A2(G257), .A3(G389), .ZN(new_n1523_));
  NOR2_X1   g1094(.A1(new_n514_), .A2(new_n568_), .ZN(new_n1524_));
  OAI21_X1  g1095(.A(new_n567_), .B1(new_n540_), .B2(G257), .ZN(new_n1525_));
  OAI211_X1 g1096(.A(new_n1522_), .B(new_n1523_), .C1(new_n1524_), .C2(new_n1525_), .ZN(new_n1526_));
  INV_X1    g1097(.A(G400), .ZN(new_n1527_));
  AOI21_X1  g1098(.A(new_n1527_), .B1(G251), .B2(new_n555_), .ZN(new_n1528_));
  OAI21_X1  g1099(.A(new_n1528_), .B1(new_n518_), .B2(new_n555_), .ZN(new_n1529_));
  NOR2_X1   g1100(.A1(new_n555_), .A2(G242), .ZN(new_n1530_));
  OAI21_X1  g1101(.A(new_n1527_), .B1(G254), .B2(G265), .ZN(new_n1531_));
  OAI21_X1  g1102(.A(new_n1529_), .B1(new_n1530_), .B2(new_n1531_), .ZN(new_n1532_));
  XNOR2_X1  g1103(.A(new_n1526_), .B(new_n1532_), .ZN(new_n1533_));
  AOI21_X1  g1104(.A(G457), .B1(G210), .B2(G242), .ZN(new_n1534_));
  INV_X1    g1105(.A(KEYINPUT120), .ZN(new_n1535_));
  AOI22_X1  g1106(.A1(new_n1534_), .A2(new_n1535_), .B1(new_n616_), .B2(G254), .ZN(new_n1536_));
  OAI21_X1  g1107(.A(new_n1536_), .B1(new_n1535_), .B2(new_n1534_), .ZN(new_n1537_));
  AOI22_X1  g1108(.A1(new_n617_), .A2(G251), .B1(G210), .B2(G248), .ZN(new_n1538_));
  OAI21_X1  g1109(.A(new_n1537_), .B1(new_n1538_), .B2(new_n620_), .ZN(new_n1539_));
  XOR2_X1   g1110(.A(new_n1533_), .B(new_n1539_), .Z(new_n1540_));
  AOI21_X1  g1111(.A(G4091), .B1(new_n1520_), .B2(new_n1540_), .ZN(new_n1541_));
  OAI21_X1  g1112(.A(new_n1541_), .B1(new_n1540_), .B2(new_n1520_), .ZN(new_n1542_));
  NOR2_X1   g1113(.A1(new_n1542_), .A2(G4092), .ZN(new_n1543_));
  XNOR2_X1  g1114(.A(new_n1543_), .B(KEYINPUT121), .ZN(new_n1544_));
  INV_X1    g1115(.A(KEYINPUT108), .ZN(new_n1545_));
  NAND2_X1  g1116(.A1(new_n945_), .A2(new_n951_), .ZN(new_n1546_));
  NAND2_X1  g1117(.A1(new_n955_), .A2(new_n956_), .ZN(new_n1547_));
  AND4_X1   g1118(.A1(new_n1545_), .A2(new_n1546_), .A3(new_n1547_), .A4(new_n961_), .ZN(new_n1548_));
  AOI21_X1  g1119(.A(new_n1545_), .B1(new_n957_), .B2(new_n961_), .ZN(new_n1549_));
  INV_X1    g1120(.A(new_n811_), .ZN(new_n1550_));
  NAND4_X1  g1121(.A1(new_n973_), .A2(new_n1550_), .A3(new_n971_), .A4(new_n972_), .ZN(new_n1551_));
  AND2_X1   g1122(.A1(new_n985_), .A2(new_n675_), .ZN(new_n1552_));
  INV_X1    g1123(.A(new_n972_), .ZN(new_n1553_));
  OAI21_X1  g1124(.A(new_n811_), .B1(new_n1552_), .B2(new_n1553_), .ZN(new_n1554_));
  AOI21_X1  g1125(.A(new_n989_), .B1(new_n1551_), .B2(new_n1554_), .ZN(new_n1555_));
  AND3_X1   g1126(.A1(new_n1551_), .A2(new_n989_), .A3(new_n1554_), .ZN(new_n1556_));
  OAI22_X1  g1127(.A1(new_n1548_), .A2(new_n1549_), .B1(new_n1555_), .B2(new_n1556_), .ZN(new_n1557_));
  NAND3_X1  g1128(.A1(new_n1546_), .A2(new_n1547_), .A3(new_n961_), .ZN(new_n1558_));
  NAND2_X1  g1129(.A1(new_n1558_), .A2(KEYINPUT108), .ZN(new_n1559_));
  NAND2_X1  g1130(.A1(new_n1551_), .A2(new_n1554_), .ZN(new_n1560_));
  AND3_X1   g1131(.A1(new_n986_), .A2(new_n987_), .A3(new_n988_), .ZN(new_n1561_));
  NAND2_X1  g1132(.A1(new_n1560_), .A2(new_n1561_), .ZN(new_n1562_));
  NAND3_X1  g1133(.A1(new_n957_), .A2(new_n1545_), .A3(new_n961_), .ZN(new_n1563_));
  NAND3_X1  g1134(.A1(new_n1551_), .A2(new_n989_), .A3(new_n1554_), .ZN(new_n1564_));
  NAND4_X1  g1135(.A1(new_n1559_), .A2(new_n1562_), .A3(new_n1563_), .A4(new_n1564_), .ZN(new_n1565_));
  AND3_X1   g1136(.A1(new_n1557_), .A2(new_n781_), .A3(new_n1565_), .ZN(new_n1566_));
  AOI21_X1  g1137(.A(new_n781_), .B1(new_n1557_), .B2(new_n1565_), .ZN(new_n1567_));
  INV_X1    g1138(.A(KEYINPUT109), .ZN(new_n1568_));
  NOR3_X1   g1139(.A1(new_n1566_), .A2(new_n1567_), .A3(new_n1568_), .ZN(new_n1569_));
  NAND2_X1  g1140(.A1(new_n1567_), .A2(new_n1568_), .ZN(new_n1570_));
  INV_X1    g1141(.A(new_n1570_), .ZN(new_n1571_));
  OAI21_X1  g1142(.A(new_n669_), .B1(new_n1569_), .B2(new_n1571_), .ZN(new_n1572_));
  INV_X1    g1143(.A(new_n669_), .ZN(new_n1573_));
  OAI21_X1  g1144(.A(new_n1573_), .B1(new_n1566_), .B2(new_n1567_), .ZN(new_n1574_));
  NAND3_X1  g1145(.A1(new_n1572_), .A2(KEYINPUT110), .A3(new_n1574_), .ZN(new_n1575_));
  INV_X1    g1146(.A(KEYINPUT110), .ZN(new_n1576_));
  OAI211_X1 g1147(.A(new_n1576_), .B(new_n669_), .C1(new_n1569_), .C2(new_n1571_), .ZN(new_n1577_));
  AOI21_X1  g1148(.A(new_n779_), .B1(new_n1575_), .B2(new_n1577_), .ZN(new_n1578_));
  AND4_X1   g1149(.A1(new_n1559_), .A2(new_n1563_), .A3(new_n1562_), .A4(new_n1564_), .ZN(new_n1579_));
  AOI22_X1  g1150(.A1(new_n1559_), .A2(new_n1563_), .B1(new_n1562_), .B2(new_n1564_), .ZN(new_n1580_));
  OAI21_X1  g1151(.A(new_n780_), .B1(new_n1579_), .B2(new_n1580_), .ZN(new_n1581_));
  NAND3_X1  g1152(.A1(new_n1557_), .A2(new_n781_), .A3(new_n1565_), .ZN(new_n1582_));
  NAND3_X1  g1153(.A1(new_n1581_), .A2(KEYINPUT109), .A3(new_n1582_), .ZN(new_n1583_));
  AOI21_X1  g1154(.A(new_n1573_), .B1(new_n1583_), .B2(new_n1570_), .ZN(new_n1584_));
  NAND2_X1  g1155(.A1(new_n1574_), .A2(KEYINPUT110), .ZN(new_n1585_));
  NOR2_X1   g1156(.A1(new_n1584_), .A2(new_n1585_), .ZN(new_n1586_));
  AOI211_X1 g1157(.A(KEYINPUT110), .B(new_n1573_), .C1(new_n1583_), .C2(new_n1570_), .ZN(new_n1587_));
  NOR3_X1   g1158(.A1(new_n1586_), .A2(new_n1587_), .A3(new_n629_), .ZN(new_n1588_));
  OAI21_X1  g1159(.A(new_n683_), .B1(new_n1578_), .B2(new_n1588_), .ZN(new_n1589_));
  AOI21_X1  g1160(.A(new_n669_), .B1(new_n1583_), .B2(new_n1570_), .ZN(new_n1590_));
  OAI21_X1  g1161(.A(new_n669_), .B1(new_n1566_), .B2(new_n1567_), .ZN(new_n1591_));
  NAND2_X1  g1162(.A1(new_n1591_), .A2(new_n779_), .ZN(new_n1592_));
  OAI21_X1  g1163(.A(new_n782_), .B1(new_n1590_), .B2(new_n1592_), .ZN(new_n1593_));
  OAI21_X1  g1164(.A(new_n1577_), .B1(new_n1584_), .B2(new_n1585_), .ZN(new_n1594_));
  AOI21_X1  g1165(.A(new_n1593_), .B1(new_n1594_), .B2(new_n629_), .ZN(new_n1595_));
  INV_X1    g1166(.A(new_n1595_), .ZN(new_n1596_));
  NAND3_X1  g1167(.A1(new_n1589_), .A2(new_n946_), .A3(new_n1596_), .ZN(new_n1597_));
  OAI21_X1  g1168(.A(new_n629_), .B1(new_n1586_), .B2(new_n1587_), .ZN(new_n1598_));
  OAI211_X1 g1169(.A(new_n1577_), .B(new_n779_), .C1(new_n1584_), .C2(new_n1585_), .ZN(new_n1599_));
  AOI21_X1  g1170(.A(new_n682_), .B1(new_n1598_), .B2(new_n1599_), .ZN(new_n1600_));
  OAI21_X1  g1171(.A(new_n643_), .B1(new_n1600_), .B2(new_n1595_), .ZN(new_n1601_));
  INV_X1    g1172(.A(G1497), .ZN(new_n1602_));
  NAND3_X1  g1173(.A1(new_n1597_), .A2(new_n1601_), .A3(new_n1602_), .ZN(new_n1603_));
  XNOR2_X1  g1174(.A(new_n705_), .B(new_n702_), .ZN(new_n1604_));
  NOR2_X1   g1175(.A1(new_n689_), .A2(new_n806_), .ZN(new_n1605_));
  INV_X1    g1176(.A(KEYINPUT99), .ZN(new_n1606_));
  AOI21_X1  g1177(.A(new_n1605_), .B1(new_n1041_), .B2(new_n1606_), .ZN(new_n1607_));
  OAI21_X1  g1178(.A(new_n1607_), .B1(new_n1606_), .B2(new_n1041_), .ZN(new_n1608_));
  XNOR2_X1  g1179(.A(new_n1044_), .B(new_n1608_), .ZN(new_n1609_));
  OR2_X1    g1180(.A1(new_n1609_), .A2(new_n694_), .ZN(new_n1610_));
  AOI21_X1  g1181(.A(new_n1604_), .B1(new_n1610_), .B2(KEYINPUT100), .ZN(new_n1611_));
  XNOR2_X1  g1182(.A(new_n1609_), .B(new_n694_), .ZN(new_n1612_));
  OR2_X1    g1183(.A1(new_n1611_), .A2(new_n1612_), .ZN(new_n1613_));
  NAND2_X1  g1184(.A1(new_n1611_), .A2(new_n1612_), .ZN(new_n1614_));
  NAND2_X1  g1185(.A1(new_n1613_), .A2(new_n1614_), .ZN(new_n1615_));
  OAI21_X1  g1186(.A(KEYINPUT101), .B1(new_n1615_), .B2(new_n712_), .ZN(new_n1616_));
  INV_X1    g1187(.A(KEYINPUT101), .ZN(new_n1617_));
  NAND4_X1  g1188(.A1(new_n1613_), .A2(new_n1617_), .A3(new_n711_), .A4(new_n1614_), .ZN(new_n1618_));
  NAND2_X1  g1189(.A1(new_n1615_), .A2(new_n712_), .ZN(new_n1619_));
  NAND2_X1  g1190(.A1(new_n685_), .A2(G1497), .ZN(new_n1620_));
  NAND2_X1  g1191(.A1(new_n1620_), .A2(new_n825_), .ZN(new_n1621_));
  NAND4_X1  g1192(.A1(new_n1616_), .A2(new_n1618_), .A3(new_n1619_), .A4(new_n1621_), .ZN(new_n1622_));
  INV_X1    g1193(.A(new_n1621_), .ZN(new_n1623_));
  INV_X1    g1194(.A(KEYINPUT106), .ZN(new_n1624_));
  NAND2_X1  g1195(.A1(new_n699_), .A2(new_n692_), .ZN(new_n1625_));
  NAND2_X1  g1196(.A1(new_n807_), .A2(new_n700_), .ZN(new_n1626_));
  NAND2_X1  g1197(.A1(new_n1625_), .A2(new_n1626_), .ZN(new_n1627_));
  NAND2_X1  g1198(.A1(new_n1627_), .A2(KEYINPUT102), .ZN(new_n1628_));
  INV_X1    g1199(.A(KEYINPUT102), .ZN(new_n1629_));
  NAND3_X1  g1200(.A1(new_n1625_), .A2(new_n1626_), .A3(new_n1629_), .ZN(new_n1630_));
  AND3_X1   g1201(.A1(new_n1628_), .A2(new_n809_), .A3(new_n1630_), .ZN(new_n1631_));
  AOI21_X1  g1202(.A(new_n809_), .B1(new_n1628_), .B2(new_n1630_), .ZN(new_n1632_));
  OAI21_X1  g1203(.A(new_n694_), .B1(new_n1631_), .B2(new_n1632_), .ZN(new_n1633_));
  NAND2_X1  g1204(.A1(new_n1628_), .A2(new_n1630_), .ZN(new_n1634_));
  INV_X1    g1205(.A(new_n809_), .ZN(new_n1635_));
  NAND2_X1  g1206(.A1(new_n1634_), .A2(new_n1635_), .ZN(new_n1636_));
  NAND3_X1  g1207(.A1(new_n1628_), .A2(new_n809_), .A3(new_n1630_), .ZN(new_n1637_));
  NAND3_X1  g1208(.A1(new_n1636_), .A2(new_n695_), .A3(new_n1637_), .ZN(new_n1638_));
  NAND3_X1  g1209(.A1(new_n1633_), .A2(new_n1638_), .A3(KEYINPUT103), .ZN(new_n1639_));
  INV_X1    g1210(.A(KEYINPUT103), .ZN(new_n1640_));
  NAND4_X1  g1211(.A1(new_n1636_), .A2(new_n1640_), .A3(new_n695_), .A4(new_n1637_), .ZN(new_n1641_));
  NAND2_X1  g1212(.A1(new_n1639_), .A2(new_n1641_), .ZN(new_n1642_));
  AOI21_X1  g1213(.A(KEYINPUT104), .B1(new_n1642_), .B2(new_n702_), .ZN(new_n1643_));
  INV_X1    g1214(.A(KEYINPUT104), .ZN(new_n1644_));
  AOI211_X1 g1215(.A(new_n1644_), .B(new_n701_), .C1(new_n1639_), .C2(new_n1641_), .ZN(new_n1645_));
  NOR2_X1   g1216(.A1(new_n1643_), .A2(new_n1645_), .ZN(new_n1646_));
  INV_X1    g1217(.A(KEYINPUT105), .ZN(new_n1647_));
  NAND3_X1  g1218(.A1(new_n1633_), .A2(new_n1638_), .A3(new_n1647_), .ZN(new_n1648_));
  AND2_X1   g1219(.A1(new_n1648_), .A2(new_n701_), .ZN(new_n1649_));
  NAND2_X1  g1220(.A1(new_n1633_), .A2(new_n1638_), .ZN(new_n1650_));
  NAND2_X1  g1221(.A1(new_n1650_), .A2(KEYINPUT105), .ZN(new_n1651_));
  NAND2_X1  g1222(.A1(new_n1649_), .A2(new_n1651_), .ZN(new_n1652_));
  NAND2_X1  g1223(.A1(new_n1652_), .A2(new_n705_), .ZN(new_n1653_));
  OAI21_X1  g1224(.A(new_n1624_), .B1(new_n1646_), .B2(new_n1653_), .ZN(new_n1654_));
  AOI21_X1  g1225(.A(new_n1045_), .B1(new_n1649_), .B2(new_n1651_), .ZN(new_n1655_));
  OAI211_X1 g1226(.A(new_n1655_), .B(KEYINPUT106), .C1(new_n1643_), .C2(new_n1645_), .ZN(new_n1656_));
  OAI22_X1  g1227(.A1(new_n1643_), .A2(new_n1645_), .B1(new_n702_), .B2(new_n1642_), .ZN(new_n1657_));
  AOI22_X1  g1228(.A1(new_n1654_), .A2(new_n1656_), .B1(new_n1045_), .B2(new_n1657_), .ZN(new_n1658_));
  OAI21_X1  g1229(.A(new_n1623_), .B1(new_n1658_), .B2(new_n712_), .ZN(new_n1659_));
  NAND2_X1  g1230(.A1(new_n1654_), .A2(new_n1656_), .ZN(new_n1660_));
  NAND2_X1  g1231(.A1(new_n1657_), .A2(new_n1045_), .ZN(new_n1661_));
  AND3_X1   g1232(.A1(new_n1660_), .A2(new_n712_), .A3(new_n1661_), .ZN(new_n1662_));
  OAI21_X1  g1233(.A(new_n1622_), .B1(new_n1659_), .B2(new_n1662_), .ZN(new_n1663_));
  AOI21_X1  g1234(.A(G374), .B1(new_n670_), .B2(new_n671_), .ZN(new_n1664_));
  OAI21_X1  g1235(.A(new_n972_), .B1(new_n1664_), .B2(new_n949_), .ZN(new_n1665_));
  NOR2_X1   g1236(.A1(new_n1664_), .A2(new_n972_), .ZN(new_n1666_));
  INV_X1    g1237(.A(new_n1666_), .ZN(new_n1667_));
  AND3_X1   g1238(.A1(new_n657_), .A2(new_n669_), .A3(new_n672_), .ZN(new_n1668_));
  OAI211_X1 g1239(.A(new_n1665_), .B(new_n1667_), .C1(new_n1668_), .C2(new_n989_), .ZN(new_n1669_));
  AOI21_X1  g1240(.A(new_n1553_), .B1(new_n657_), .B2(new_n783_), .ZN(new_n1670_));
  OAI211_X1 g1241(.A(new_n673_), .B(new_n1561_), .C1(new_n1670_), .C2(new_n1666_), .ZN(new_n1671_));
  INV_X1    g1242(.A(KEYINPUT107), .ZN(new_n1672_));
  NAND3_X1  g1243(.A1(new_n1669_), .A2(new_n1671_), .A3(new_n1672_), .ZN(new_n1673_));
  INV_X1    g1244(.A(new_n1558_), .ZN(new_n1674_));
  NAND2_X1  g1245(.A1(new_n1561_), .A2(new_n673_), .ZN(new_n1675_));
  NAND4_X1  g1246(.A1(new_n1675_), .A2(KEYINPUT107), .A3(new_n1665_), .A4(new_n1667_), .ZN(new_n1676_));
  NAND4_X1  g1247(.A1(new_n1673_), .A2(new_n1674_), .A3(new_n785_), .A4(new_n1676_), .ZN(new_n1677_));
  NAND3_X1  g1248(.A1(new_n957_), .A2(new_n785_), .A3(new_n961_), .ZN(new_n1678_));
  NAND3_X1  g1249(.A1(new_n1678_), .A2(new_n1669_), .A3(new_n1671_), .ZN(new_n1679_));
  AND3_X1   g1250(.A1(new_n1677_), .A2(new_n781_), .A3(new_n1679_), .ZN(new_n1680_));
  AOI21_X1  g1251(.A(new_n781_), .B1(new_n1677_), .B2(new_n1679_), .ZN(new_n1681_));
  OAI21_X1  g1252(.A(new_n1573_), .B1(new_n1680_), .B2(new_n1681_), .ZN(new_n1682_));
  NAND3_X1  g1253(.A1(new_n1677_), .A2(new_n781_), .A3(new_n1679_), .ZN(new_n1683_));
  NAND3_X1  g1254(.A1(new_n1673_), .A2(new_n1678_), .A3(new_n1676_), .ZN(new_n1684_));
  NAND3_X1  g1255(.A1(new_n1674_), .A2(new_n1669_), .A3(new_n1671_), .ZN(new_n1685_));
  NAND3_X1  g1256(.A1(new_n1684_), .A2(new_n1685_), .A3(new_n780_), .ZN(new_n1686_));
  NAND3_X1  g1257(.A1(new_n1683_), .A2(new_n669_), .A3(new_n1686_), .ZN(new_n1687_));
  AND3_X1   g1258(.A1(new_n1682_), .A2(new_n629_), .A3(new_n1687_), .ZN(new_n1688_));
  AOI21_X1  g1259(.A(new_n629_), .B1(new_n1682_), .B2(new_n1687_), .ZN(new_n1689_));
  OAI21_X1  g1260(.A(new_n683_), .B1(new_n1688_), .B2(new_n1689_), .ZN(new_n1690_));
  NAND3_X1  g1261(.A1(new_n1682_), .A2(new_n629_), .A3(new_n1687_), .ZN(new_n1691_));
  OAI21_X1  g1262(.A(new_n669_), .B1(new_n1680_), .B2(new_n1681_), .ZN(new_n1692_));
  NAND3_X1  g1263(.A1(new_n1683_), .A2(new_n1573_), .A3(new_n1686_), .ZN(new_n1693_));
  NAND3_X1  g1264(.A1(new_n1692_), .A2(new_n779_), .A3(new_n1693_), .ZN(new_n1694_));
  NAND3_X1  g1265(.A1(new_n1691_), .A2(new_n1694_), .A3(new_n782_), .ZN(new_n1695_));
  NAND3_X1  g1266(.A1(new_n1690_), .A2(new_n946_), .A3(new_n1695_), .ZN(new_n1696_));
  NAND2_X1  g1267(.A1(new_n1696_), .A2(KEYINPUT112), .ZN(new_n1697_));
  INV_X1    g1268(.A(KEYINPUT112), .ZN(new_n1698_));
  NAND4_X1  g1269(.A1(new_n1690_), .A2(new_n1698_), .A3(new_n946_), .A4(new_n1695_), .ZN(new_n1699_));
  NAND2_X1  g1270(.A1(new_n1690_), .A2(new_n1695_), .ZN(new_n1700_));
  NAND2_X1  g1271(.A1(new_n1700_), .A2(new_n643_), .ZN(new_n1701_));
  NAND3_X1  g1272(.A1(new_n1697_), .A2(new_n1699_), .A3(new_n1701_), .ZN(new_n1702_));
  AOI21_X1  g1273(.A(new_n1663_), .B1(new_n1702_), .B2(G1497), .ZN(new_n1703_));
  NAND2_X1  g1274(.A1(new_n1603_), .A2(new_n1703_), .ZN(new_n1704_));
  INV_X1    g1275(.A(KEYINPUT113), .ZN(new_n1705_));
  NAND2_X1  g1276(.A1(new_n1704_), .A2(new_n1705_), .ZN(new_n1706_));
  NAND3_X1  g1277(.A1(new_n1603_), .A2(new_n1703_), .A3(KEYINPUT113), .ZN(new_n1707_));
  NAND2_X1  g1278(.A1(new_n1706_), .A2(new_n1707_), .ZN(new_n1708_));
  INV_X1    g1279(.A(new_n1663_), .ZN(new_n1709_));
  NAND2_X1  g1280(.A1(new_n1597_), .A2(KEYINPUT111), .ZN(new_n1710_));
  INV_X1    g1281(.A(KEYINPUT111), .ZN(new_n1711_));
  NAND4_X1  g1282(.A1(new_n1589_), .A2(new_n1596_), .A3(new_n1711_), .A4(new_n946_), .ZN(new_n1712_));
  NAND4_X1  g1283(.A1(new_n1710_), .A2(new_n1602_), .A3(new_n1712_), .A4(new_n1601_), .ZN(new_n1713_));
  OR3_X1    g1284(.A1(new_n1688_), .A2(new_n1689_), .A3(new_n683_), .ZN(new_n1714_));
  NAND2_X1  g1285(.A1(new_n1691_), .A2(new_n1694_), .ZN(new_n1715_));
  NAND2_X1  g1286(.A1(new_n1715_), .A2(new_n948_), .ZN(new_n1716_));
  AOI21_X1  g1287(.A(new_n644_), .B1(new_n1714_), .B2(new_n1716_), .ZN(new_n1717_));
  INV_X1    g1288(.A(new_n1696_), .ZN(new_n1718_));
  OAI21_X1  g1289(.A(G1497), .B1(new_n1717_), .B2(new_n1718_), .ZN(new_n1719_));
  AOI21_X1  g1290(.A(new_n1709_), .B1(new_n1713_), .B2(new_n1719_), .ZN(new_n1720_));
  OAI21_X1  g1291(.A(G4091), .B1(new_n1708_), .B2(new_n1720_), .ZN(new_n1721_));
  OAI211_X1 g1292(.A(new_n1487_), .B(new_n1544_), .C1(new_n1721_), .C2(G4092), .ZN(G882));
  OAI21_X1  g1293(.A(G4087), .B1(G14), .B2(G4088), .ZN(new_n1723_));
  INV_X1    g1294(.A(G64), .ZN(new_n1724_));
  AOI21_X1  g1295(.A(new_n1723_), .B1(new_n1724_), .B2(G4088), .ZN(new_n1725_));
  INV_X1    g1296(.A(KEYINPUT124), .ZN(new_n1726_));
  NAND2_X1  g1297(.A1(G94), .A2(G4092), .ZN(new_n1727_));
  OR2_X1    g1298(.A1(new_n1727_), .A2(KEYINPUT123), .ZN(new_n1728_));
  NAND2_X1  g1299(.A1(new_n1727_), .A2(KEYINPUT123), .ZN(new_n1729_));
  NAND2_X1  g1300(.A1(new_n1728_), .A2(new_n1729_), .ZN(new_n1730_));
  AND3_X1   g1301(.A1(new_n1481_), .A2(new_n1388_), .A3(new_n1482_), .ZN(new_n1731_));
  AOI21_X1  g1302(.A(new_n1482_), .B1(new_n1481_), .B2(new_n1388_), .ZN(new_n1732_));
  OAI21_X1  g1303(.A(G4091), .B1(new_n1731_), .B2(new_n1732_), .ZN(new_n1733_));
  AOI21_X1  g1304(.A(G4092), .B1(new_n1365_), .B2(new_n855_), .ZN(new_n1734_));
  AOI21_X1  g1305(.A(new_n1730_), .B1(new_n1733_), .B2(new_n1734_), .ZN(new_n1735_));
  OAI21_X1  g1306(.A(new_n1726_), .B1(new_n1735_), .B2(new_n1097_), .ZN(new_n1736_));
  INV_X1    g1307(.A(new_n1734_), .ZN(new_n1737_));
  AOI21_X1  g1308(.A(new_n1737_), .B1(new_n1484_), .B2(G4091), .ZN(new_n1738_));
  OAI211_X1 g1309(.A(KEYINPUT124), .B(new_n1096_), .C1(new_n1738_), .C2(new_n1730_), .ZN(new_n1739_));
  AOI21_X1  g1310(.A(new_n1725_), .B1(new_n1736_), .B2(new_n1739_), .ZN(new_n1740_));
  NAND2_X1  g1311(.A1(new_n1542_), .A2(new_n847_), .ZN(new_n1741_));
  INV_X1    g1312(.A(new_n1741_), .ZN(new_n1742_));
  AOI22_X1  g1313(.A1(new_n1721_), .A2(new_n1742_), .B1(G97), .B2(G4092), .ZN(new_n1743_));
  INV_X1    g1314(.A(KEYINPUT122), .ZN(new_n1744_));
  NOR3_X1   g1315(.A1(new_n1743_), .A2(new_n1744_), .A3(new_n902_), .ZN(new_n1745_));
  NAND2_X1  g1316(.A1(G97), .A2(G4092), .ZN(new_n1746_));
  AND3_X1   g1317(.A1(new_n1603_), .A2(new_n1703_), .A3(KEYINPUT113), .ZN(new_n1747_));
  AOI21_X1  g1318(.A(KEYINPUT113), .B1(new_n1603_), .B2(new_n1703_), .ZN(new_n1748_));
  NOR2_X1   g1319(.A1(new_n1747_), .A2(new_n1748_), .ZN(new_n1749_));
  NOR3_X1   g1320(.A1(new_n1600_), .A2(new_n643_), .A3(new_n1595_), .ZN(new_n1750_));
  OAI211_X1 g1321(.A(new_n1602_), .B(new_n1601_), .C1(new_n1750_), .C2(new_n1711_), .ZN(new_n1751_));
  INV_X1    g1322(.A(new_n1712_), .ZN(new_n1752_));
  OAI21_X1  g1323(.A(new_n1719_), .B1(new_n1751_), .B2(new_n1752_), .ZN(new_n1753_));
  NAND2_X1  g1324(.A1(new_n1753_), .A2(new_n1663_), .ZN(new_n1754_));
  AOI21_X1  g1325(.A(new_n855_), .B1(new_n1749_), .B2(new_n1754_), .ZN(new_n1755_));
  OAI21_X1  g1326(.A(new_n1746_), .B1(new_n1755_), .B2(new_n1741_), .ZN(new_n1756_));
  AOI21_X1  g1327(.A(KEYINPUT122), .B1(new_n1756_), .B2(new_n901_), .ZN(new_n1757_));
  OAI21_X1  g1328(.A(new_n1740_), .B1(new_n1745_), .B2(new_n1757_), .ZN(G767));
  NAND2_X1  g1329(.A1(new_n1724_), .A2(G4089), .ZN(new_n1759_));
  OAI211_X1 g1330(.A(new_n1759_), .B(G4090), .C1(G14), .C2(G4089), .ZN(new_n1760_));
  AOI21_X1  g1331(.A(new_n855_), .B1(new_n1478_), .B2(new_n1483_), .ZN(new_n1761_));
  OAI211_X1 g1332(.A(new_n1729_), .B(new_n1728_), .C1(new_n1761_), .C2(new_n1737_), .ZN(new_n1762_));
  AOI21_X1  g1333(.A(KEYINPUT125), .B1(new_n1762_), .B2(new_n1112_), .ZN(new_n1763_));
  INV_X1    g1334(.A(KEYINPUT125), .ZN(new_n1764_));
  NOR3_X1   g1335(.A1(new_n1735_), .A2(new_n1764_), .A3(new_n1124_), .ZN(new_n1765_));
  OAI221_X1 g1336(.A(new_n1760_), .B1(new_n940_), .B2(new_n1743_), .C1(new_n1763_), .C2(new_n1765_), .ZN(G807));
  NAND3_X1  g1337(.A1(new_n1071_), .A2(G176), .A3(G1690), .ZN(new_n1767_));
  OR2_X1    g1338(.A1(new_n1767_), .A2(KEYINPUT126), .ZN(new_n1768_));
  NAND3_X1  g1339(.A1(G179), .A2(G1689), .A3(G1690), .ZN(new_n1769_));
  NAND2_X1  g1340(.A1(new_n1767_), .A2(KEYINPUT126), .ZN(new_n1770_));
  NAND3_X1  g1341(.A1(new_n1768_), .A2(new_n1769_), .A3(new_n1770_), .ZN(new_n1771_));
  AOI21_X1  g1342(.A(new_n1771_), .B1(new_n1762_), .B2(new_n1078_), .ZN(new_n1772_));
  INV_X1    g1343(.A(new_n1072_), .ZN(new_n1773_));
  OAI21_X1  g1344(.A(new_n1772_), .B1(new_n1773_), .B2(new_n1743_), .ZN(new_n1774_));
  NAND2_X1  g1345(.A1(new_n1774_), .A2(G137), .ZN(G658));
  NAND3_X1  g1346(.A1(new_n1081_), .A2(G176), .A3(G1694), .ZN(new_n1776_));
  INV_X1    g1347(.A(KEYINPUT127), .ZN(new_n1777_));
  OR2_X1    g1348(.A1(new_n1776_), .A2(new_n1777_), .ZN(new_n1778_));
  NAND3_X1  g1349(.A1(G179), .A2(G1691), .A3(G1694), .ZN(new_n1779_));
  NAND2_X1  g1350(.A1(new_n1776_), .A2(new_n1777_), .ZN(new_n1780_));
  NAND3_X1  g1351(.A1(new_n1778_), .A2(new_n1779_), .A3(new_n1780_), .ZN(new_n1781_));
  AOI21_X1  g1352(.A(new_n1781_), .B1(new_n1762_), .B2(new_n1167_), .ZN(new_n1782_));
  OAI21_X1  g1353(.A(new_n1782_), .B1(new_n1083_), .B2(new_n1743_), .ZN(new_n1783_));
  NAND2_X1  g1354(.A1(new_n1783_), .A2(G137), .ZN(G690));
endmodule


