//Secret key is'1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_c7552" written by ABC on Wed Nov  2 14:11:17 2022

module locked_c7552 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G5, G9, G12, G15,
    G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55,
    G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87,
    G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113,
    G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141,
    G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159,
    G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171,
    G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183,
    G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195,
    G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207,
    G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219,
    G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231,
    G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197,
    G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208,
    G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698,
    G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393,
    G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526,
    G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G5, G9,
    G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53,
    G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69,
    G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85,
    G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112,
    G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138,
    G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158,
    G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170,
    G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218,
    G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230,
    G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339,
    G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204,
    G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256,
    G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749,
    G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437,
    G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_n426_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1102_, new_n1103_,
    new_n1105_, new_n1106_, new_n1108_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1271_,
    new_n1272_, new_n1273_, new_n1276_, new_n1277_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1304_, new_n1305_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1326_, new_n1327_, new_n1328_, new_n1331_, new_n1332_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1347_, new_n1350_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1380_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1400_, new_n1401_, new_n1402_,
    new_n1404_, new_n1406_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_;
  BUF_X1    g0000(.A(G1), .Z(G2));
  BUF_X1    g0001(.A(G1), .Z(G3));
  BUF_X1    g0002(.A(G1459), .Z(G450));
  BUF_X1    g0003(.A(G1469), .Z(G448));
  BUF_X1    g0004(.A(G1480), .Z(G444));
  BUF_X1    g0005(.A(G1486), .Z(G442));
  BUF_X1    g0006(.A(G1492), .Z(G440));
  BUF_X1    g0007(.A(G1496), .Z(G438));
  BUF_X1    g0008(.A(G2208), .Z(G496));
  BUF_X1    g0009(.A(G2218), .Z(G494));
  BUF_X1    g0010(.A(G2224), .Z(G492));
  XNOR2_X1  g0011(.A(KEYINPUT0), .B(G2230), .ZN(G490));
  BUF_X1    g0012(.A(G2236), .Z(G488));
  BUF_X1    g0013(.A(G2239), .Z(G486));
  BUF_X1    g0014(.A(G2247), .Z(G484));
  BUF_X1    g0015(.A(G2253), .Z(G482));
  BUF_X1    g0016(.A(G2256), .Z(G480));
  BUF_X1    g0017(.A(G3698), .Z(G560));
  BUF_X1    g0018(.A(G3701), .Z(G542));
  BUF_X1    g0019(.A(G3705), .Z(G558));
  BUF_X1    g0020(.A(G3711), .Z(G556));
  BUF_X1    g0021(.A(G3717), .Z(G554));
  BUF_X1    g0022(.A(G3723), .Z(G552));
  BUF_X1    g0023(.A(G3729), .Z(G550));
  BUF_X1    g0024(.A(G3737), .Z(G548));
  BUF_X1    g0025(.A(G3743), .Z(G546));
  BUF_X1    g0026(.A(G3749), .Z(G544));
  BUF_X1    g0027(.A(G4393), .Z(G540));
  XNOR2_X1  g0028(.A(KEYINPUT1), .B(G4400), .ZN(G538));
  BUF_X1    g0029(.A(G4405), .Z(G536));
  BUF_X1    g0030(.A(G4410), .Z(G534));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G4415), .Z(G532));
  BUF_X1    g0032(.A(G4420), .Z(G530));
  BUF_X1    g0033(.A(G4427), .Z(G528));
  BUF_X1    g0034(.A(G4432), .Z(G526));
  BUF_X1    g0035(.A(G4437), .Z(G524));
  INV_X1    g0036(.A(G15), .ZN(G279));
  BUF_X1    g0037(.A(G1462), .Z(G436));
  BUF_X1    g0038(.A(G2211), .Z(G478));
  BUF_X1    g0039(.A(G4394), .Z(G522));
  OR2_X1    g0040(.A1(G5), .A2(G57), .ZN(G402));
  NAND4_X1  g0041(.A1(G150), .A2(G184), .A3(G228), .A4(G240), .ZN(G404));
  NAND4_X1  g0042(.A1(G152), .A2(G210), .A3(G218), .A4(G230), .ZN(G406));
  NAND4_X1  g0043(.A1(G182), .A2(G183), .A3(G185), .A4(G186), .ZN(G408));
  NAND4_X1  g0044(.A1(G162), .A2(G172), .A3(G188), .A4(G199), .ZN(G410));
  BUF_X1    g0045(.A(G1), .Z(G432));
  BUF_X1    g0046(.A(G106), .Z(G446));
  INV_X1    g0047(.A(G5), .ZN(new_n426_));
  NAND2_X1  g0048(.A1(new_n426_), .A2(G1197), .ZN(G284));
  INV_X1    g0049(.A(G15), .ZN(G286));
  NAND2_X1  g0050(.A1(new_n426_), .A2(G1197), .ZN(G289));
  NAND3_X1  g0051(.A1(new_n426_), .A2(G133), .A3(G134), .ZN(G292));
  INV_X1    g0052(.A(G15), .ZN(G341));
  NAND3_X1  g0053(.A1(new_n426_), .A2(G133), .A3(G134), .ZN(G281));
  BUF_X1    g0054(.A(G1), .Z(G453));
  AND2_X1   g0055(.A1(G1), .A2(G163), .ZN(G278));
  INV_X1    g0056(.A(G41), .ZN(new_n435_));
  NOR3_X1   g0057(.A1(new_n435_), .A2(G18), .A3(G3701), .ZN(new_n436_));
  INV_X1    g0058(.A(G3701), .ZN(new_n437_));
  NOR3_X1   g0059(.A1(new_n437_), .A2(G18), .A3(G41), .ZN(new_n438_));
  NOR2_X1   g0060(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g0061(.A(G4526), .ZN(new_n440_));
  XNOR2_X1  g0062(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g0063(.A(new_n441_), .B(KEYINPUT3), .ZN(G373));
  INV_X1    g0064(.A(G154), .ZN(new_n443_));
  NAND2_X1  g0065(.A1(new_n443_), .A2(KEYINPUT5), .ZN(new_n444_));
  INV_X1    g0066(.A(KEYINPUT5), .ZN(new_n445_));
  NAND2_X1  g0067(.A1(new_n445_), .A2(G154), .ZN(new_n446_));
  NAND3_X1  g0068(.A1(new_n444_), .A2(new_n446_), .A3(G18), .ZN(new_n447_));
  NAND2_X1  g0069(.A1(G9), .A2(G12), .ZN(new_n448_));
  NAND2_X1  g0070(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g0071(.A1(new_n449_), .A2(G2253), .ZN(new_n450_));
  INV_X1    g0072(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g0073(.A1(new_n449_), .A2(G2253), .ZN(new_n452_));
  NAND2_X1  g0074(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g0075(.A(new_n448_), .ZN(new_n454_));
  INV_X1    g0076(.A(G156), .ZN(new_n455_));
  AOI21_X1  g0077(.A(new_n454_), .B1(G18), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g0078(.A(G2239), .ZN(new_n457_));
  NAND2_X1  g0079(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g0080(.A(G155), .ZN(new_n459_));
  AOI21_X1  g0081(.A(new_n454_), .B1(G18), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g0082(.A(G2247), .ZN(new_n461_));
  NAND2_X1  g0083(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g0084(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g0085(.A(new_n463_), .B1(new_n461_), .B2(new_n460_), .ZN(new_n464_));
  NOR2_X1   g0086(.A1(new_n453_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g0087(.A1(new_n465_), .A2(new_n450_), .ZN(new_n466_));
  INV_X1    g0088(.A(G18), .ZN(new_n467_));
  OAI21_X1  g0089(.A(new_n448_), .B1(new_n467_), .B2(G153), .ZN(new_n468_));
  XNOR2_X1  g0090(.A(new_n468_), .B(KEYINPUT6), .ZN(new_n469_));
  AND2_X1   g0091(.A1(new_n469_), .A2(G2256), .ZN(new_n470_));
  NOR2_X1   g0092(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g0093(.A1(new_n469_), .A2(G2256), .ZN(new_n472_));
  INV_X1    g0094(.A(G135), .ZN(new_n473_));
  NOR2_X1   g0095(.A1(new_n473_), .A2(G18), .ZN(new_n474_));
  AOI21_X1  g0096(.A(new_n474_), .B1(G18), .B2(G158), .ZN(new_n475_));
  OR2_X1    g0097(.A1(new_n475_), .A2(G2230), .ZN(new_n476_));
  INV_X1    g0098(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g0099(.A1(new_n467_), .A2(G138), .ZN(new_n478_));
  NAND2_X1  g0100(.A1(G18), .A2(G160), .ZN(new_n479_));
  AND2_X1   g0101(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g0102(.A(G2218), .ZN(new_n481_));
  AOI21_X1  g0103(.A(new_n480_), .B1(KEYINPUT9), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g0104(.A(new_n482_), .B1(KEYINPUT9), .B2(new_n481_), .ZN(new_n483_));
  INV_X1    g0105(.A(new_n480_), .ZN(new_n484_));
  OR3_X1    g0106(.A1(new_n484_), .A2(KEYINPUT9), .A3(new_n481_), .ZN(new_n485_));
  NAND2_X1  g0107(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g0108(.A(KEYINPUT8), .B(G144), .Z(new_n487_));
  NAND2_X1  g0109(.A1(new_n487_), .A2(new_n467_), .ZN(new_n488_));
  NAND2_X1  g0110(.A1(G18), .A2(G159), .ZN(new_n489_));
  NAND2_X1  g0111(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g0112(.A(G2224), .ZN(new_n491_));
  NAND2_X1  g0113(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g0114(.A1(new_n489_), .A2(G2224), .ZN(new_n493_));
  INV_X1    g0115(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g0116(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g0117(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g0118(.A1(new_n486_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g0119(.A1(new_n467_), .A2(G147), .ZN(new_n498_));
  AOI21_X1  g0120(.A(new_n498_), .B1(G18), .B2(G151), .ZN(new_n499_));
  OR2_X1    g0121(.A1(new_n499_), .A2(G2211), .ZN(new_n500_));
  INV_X1    g0122(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g0123(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g0124(.A1(new_n502_), .A2(new_n492_), .ZN(new_n503_));
  NAND2_X1  g0125(.A1(new_n475_), .A2(G2230), .ZN(new_n504_));
  AOI21_X1  g0126(.A(new_n477_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g0127(.A(new_n448_), .B1(new_n467_), .B2(G157), .ZN(new_n506_));
  XNOR2_X1  g0128(.A(new_n506_), .B(KEYINPUT7), .ZN(new_n507_));
  INV_X1    g0129(.A(G2236), .ZN(new_n508_));
  NAND2_X1  g0130(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g0131(.A1(new_n476_), .A2(new_n504_), .ZN(new_n510_));
  NOR2_X1   g0132(.A1(new_n496_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g0133(.A1(new_n484_), .A2(new_n481_), .ZN(new_n512_));
  INV_X1    g0134(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g0135(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g0136(.A1(new_n505_), .A2(new_n509_), .A3(new_n514_), .ZN(new_n515_));
  OR2_X1    g0137(.A1(new_n507_), .A2(new_n508_), .ZN(new_n516_));
  AND2_X1   g0138(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g0139(.A1(new_n456_), .A2(new_n457_), .ZN(new_n518_));
  NAND2_X1  g0140(.A1(new_n518_), .A2(new_n462_), .ZN(new_n519_));
  NOR2_X1   g0141(.A1(new_n460_), .A2(new_n461_), .ZN(new_n520_));
  OAI21_X1  g0142(.A(new_n519_), .B1(new_n520_), .B2(new_n518_), .ZN(new_n521_));
  XNOR2_X1  g0143(.A(new_n521_), .B(new_n453_), .ZN(new_n522_));
  NOR2_X1   g0144(.A1(new_n520_), .A2(new_n518_), .ZN(new_n523_));
  NAND3_X1  g0145(.A1(new_n523_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n524_));
  INV_X1    g0146(.A(new_n462_), .ZN(new_n525_));
  NOR2_X1   g0147(.A1(new_n525_), .A2(new_n520_), .ZN(new_n526_));
  INV_X1    g0148(.A(new_n458_), .ZN(new_n527_));
  NOR2_X1   g0149(.A1(new_n527_), .A2(new_n518_), .ZN(new_n528_));
  OAI21_X1  g0150(.A(new_n524_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g0151(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g0152(.A(new_n522_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g0153(.A(new_n524_), .ZN(new_n532_));
  OAI211_X1 g0154(.A(new_n451_), .B(new_n452_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n533_));
  NAND2_X1  g0155(.A1(new_n533_), .A2(new_n451_), .ZN(new_n534_));
  OR2_X1    g0156(.A1(new_n470_), .A2(new_n472_), .ZN(new_n535_));
  XOR2_X1   g0157(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  NAND3_X1  g0158(.A1(new_n531_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g0159(.A(new_n537_), .ZN(new_n538_));
  AOI211_X1 g0160(.A(new_n471_), .B(new_n472_), .C1(new_n517_), .C2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g0161(.A1(new_n499_), .A2(G2211), .ZN(new_n540_));
  NAND2_X1  g0162(.A1(new_n500_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g0163(.A1(new_n486_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g0164(.A1(new_n542_), .A2(new_n511_), .ZN(new_n543_));
  NAND2_X1  g0165(.A1(new_n516_), .A2(new_n509_), .ZN(new_n544_));
  NOR2_X1   g0166(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g0167(.A(new_n545_), .B(KEYINPUT10), .ZN(new_n546_));
  NAND2_X1  g0168(.A1(new_n538_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g0169(.A(G4427), .ZN(new_n548_));
  NOR2_X1   g0170(.A1(new_n548_), .A2(KEYINPUT16), .ZN(new_n549_));
  INV_X1    g0171(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n551_));
  NAND2_X1  g0173(.A1(new_n467_), .A2(G32), .ZN(new_n552_));
  NAND2_X1  g0174(.A1(G18), .A2(G221), .ZN(new_n553_));
  NAND2_X1  g0175(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g0176(.A(KEYINPUT15), .ZN(new_n555_));
  NAND2_X1  g0177(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g0178(.A1(new_n552_), .A2(KEYINPUT15), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g0179(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n559_));
  NOR2_X1   g0181(.A1(new_n559_), .A2(G4427), .ZN(new_n560_));
  INV_X1    g0182(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g0183(.A(new_n551_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  AOI211_X1 g0184(.A(KEYINPUT17), .B(new_n560_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n563_));
  OAI21_X1  g0185(.A(new_n550_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g0186(.A(new_n557_), .ZN(new_n565_));
  AOI21_X1  g0187(.A(KEYINPUT15), .B1(new_n552_), .B2(new_n553_), .ZN(new_n566_));
  NOR2_X1   g0188(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g0189(.A(KEYINPUT17), .B1(new_n567_), .B2(new_n560_), .ZN(new_n568_));
  NAND3_X1  g0190(.A1(new_n558_), .A2(new_n551_), .A3(new_n561_), .ZN(new_n569_));
  NAND3_X1  g0191(.A1(new_n568_), .A2(new_n549_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g0192(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g0193(.A1(new_n467_), .A2(G35), .ZN(new_n572_));
  AOI21_X1  g0194(.A(new_n572_), .B1(G18), .B2(G222), .ZN(new_n573_));
  NAND2_X1  g0195(.A1(new_n573_), .A2(G4420), .ZN(new_n574_));
  INV_X1    g0196(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g0197(.A1(new_n573_), .A2(G4420), .ZN(new_n576_));
  NOR2_X1   g0198(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g0199(.A1(new_n467_), .A2(G66), .ZN(new_n578_));
  INV_X1    g0200(.A(G219), .ZN(new_n579_));
  OAI21_X1  g0201(.A(new_n578_), .B1(new_n467_), .B2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g0202(.A(new_n580_), .B(G4437), .ZN(new_n581_));
  NAND2_X1  g0203(.A1(new_n467_), .A2(G50), .ZN(new_n582_));
  INV_X1    g0204(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g0205(.A(new_n583_), .B1(G18), .B2(G220), .ZN(new_n584_));
  NAND2_X1  g0206(.A1(new_n584_), .A2(G4432), .ZN(new_n585_));
  INV_X1    g0207(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g0208(.A1(new_n584_), .A2(G4432), .ZN(new_n587_));
  NOR2_X1   g0209(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g0210(.A1(new_n571_), .A2(new_n577_), .A3(new_n581_), .A4(new_n588_), .ZN(new_n589_));
  INV_X1    g0211(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g0212(.A1(new_n467_), .A2(G47), .ZN(new_n591_));
  NAND2_X1  g0213(.A1(G18), .A2(G223), .ZN(new_n592_));
  AND2_X1   g0214(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OR2_X1    g0215(.A1(new_n593_), .A2(G4415), .ZN(new_n594_));
  NAND2_X1  g0216(.A1(new_n593_), .A2(G4415), .ZN(new_n595_));
  NAND2_X1  g0217(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g0218(.A1(new_n467_), .A2(G94), .ZN(new_n597_));
  NAND2_X1  g0219(.A1(G18), .A2(G225), .ZN(new_n598_));
  NAND2_X1  g0220(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g0221(.A(G4405), .ZN(new_n600_));
  NAND2_X1  g0222(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g0223(.A1(new_n597_), .A2(G4405), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g0224(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g0225(.A1(new_n596_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g0226(.A1(new_n467_), .A2(G121), .ZN(new_n605_));
  AOI21_X1  g0227(.A(new_n605_), .B1(G18), .B2(G224), .ZN(new_n606_));
  NAND2_X1  g0228(.A1(new_n606_), .A2(G4410), .ZN(new_n607_));
  INV_X1    g0229(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g0230(.A1(new_n606_), .A2(G4410), .ZN(new_n609_));
  NOR2_X1   g0231(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g0232(.A1(new_n467_), .A2(G97), .ZN(new_n611_));
  NAND2_X1  g0233(.A1(G18), .A2(G226), .ZN(new_n612_));
  NAND3_X1  g0234(.A1(new_n611_), .A2(G4400), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g0235(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g0236(.A(G4400), .B1(new_n611_), .B2(new_n612_), .ZN(new_n615_));
  NOR2_X1   g0237(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g0238(.A1(new_n467_), .A2(G118), .ZN(new_n617_));
  INV_X1    g0239(.A(G217), .ZN(new_n618_));
  OAI21_X1  g0240(.A(new_n617_), .B1(new_n467_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g0241(.A(G4394), .ZN(new_n620_));
  NAND2_X1  g0242(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g0243(.A(new_n617_), .B(G4394), .C1(new_n467_), .C2(new_n618_), .ZN(new_n622_));
  NAND2_X1  g0244(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g0245(.A(new_n623_), .ZN(new_n624_));
  NAND4_X1  g0246(.A1(new_n604_), .A2(new_n610_), .A3(new_n616_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g0247(.A(new_n625_), .ZN(new_n626_));
  AND2_X1   g0248(.A1(G18), .A2(G231), .ZN(new_n627_));
  AOI21_X1  g0249(.A(new_n627_), .B1(new_n467_), .B2(G100), .ZN(new_n628_));
  NAND2_X1  g0250(.A1(new_n628_), .A2(G3749), .ZN(new_n629_));
  INV_X1    g0251(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g0252(.A(KEYINPUT12), .ZN(new_n631_));
  OR2_X1    g0253(.A1(new_n631_), .A2(G235), .ZN(new_n632_));
  NAND2_X1  g0254(.A1(new_n631_), .A2(G235), .ZN(new_n633_));
  NAND3_X1  g0255(.A1(new_n632_), .A2(new_n633_), .A3(G18), .ZN(new_n634_));
  NAND2_X1  g0256(.A1(new_n467_), .A2(G103), .ZN(new_n635_));
  NAND2_X1  g0257(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g0258(.A(G3723), .ZN(new_n637_));
  NAND2_X1  g0259(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g0260(.A(KEYINPUT11), .B(G3711), .ZN(new_n639_));
  NAND2_X1  g0261(.A1(new_n467_), .A2(G26), .ZN(new_n640_));
  NAND2_X1  g0262(.A1(G18), .A2(G237), .ZN(new_n641_));
  NAND2_X1  g0263(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g0264(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g0265(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g0266(.A(new_n642_), .ZN(new_n645_));
  OAI21_X1  g0267(.A(new_n644_), .B1(G3711), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g0268(.A1(G18), .A2(G236), .ZN(new_n647_));
  INV_X1    g0269(.A(G23), .ZN(new_n648_));
  OAI21_X1  g0270(.A(new_n647_), .B1(new_n648_), .B2(G18), .ZN(new_n649_));
  INV_X1    g0271(.A(new_n649_), .ZN(new_n650_));
  OR2_X1    g0272(.A1(new_n650_), .A2(G3717), .ZN(new_n651_));
  NAND2_X1  g0273(.A1(new_n650_), .A2(G3717), .ZN(new_n652_));
  NAND2_X1  g0274(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g0275(.A(G29), .ZN(new_n654_));
  INV_X1    g0276(.A(G238), .ZN(new_n655_));
  MUX2_X1   g0277(.A(new_n654_), .B(new_n655_), .S(G18), .Z(new_n656_));
  NAND2_X1  g0278(.A1(new_n656_), .A2(G3705), .ZN(new_n657_));
  NAND2_X1  g0279(.A1(new_n467_), .A2(G29), .ZN(new_n658_));
  OAI21_X1  g0280(.A(new_n658_), .B1(new_n467_), .B2(new_n655_), .ZN(new_n659_));
  INV_X1    g0281(.A(G3705), .ZN(new_n660_));
  NAND2_X1  g0282(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0283(.A1(new_n657_), .A2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g0284(.A1(new_n646_), .A2(new_n653_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g0285(.A(new_n636_), .B(G3723), .ZN(new_n664_));
  NAND4_X1  g0286(.A1(new_n663_), .A2(G4526), .A3(new_n439_), .A4(new_n664_), .ZN(new_n665_));
  INV_X1    g0287(.A(new_n651_), .ZN(new_n666_));
  NAND2_X1  g0288(.A1(new_n639_), .A2(new_n642_), .ZN(new_n667_));
  INV_X1    g0289(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g0290(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g0291(.A(new_n661_), .ZN(new_n670_));
  AOI21_X1  g0292(.A(new_n670_), .B1(new_n436_), .B2(new_n657_), .ZN(new_n671_));
  OAI21_X1  g0293(.A(new_n669_), .B1(new_n671_), .B2(new_n646_), .ZN(new_n672_));
  AOI21_X1  g0294(.A(new_n666_), .B1(new_n672_), .B2(new_n652_), .ZN(new_n673_));
  NOR2_X1   g0295(.A1(new_n636_), .A2(new_n637_), .ZN(new_n674_));
  OAI211_X1 g0296(.A(new_n638_), .B(new_n665_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n675_));
  AND2_X1   g0297(.A1(G18), .A2(G232), .ZN(new_n676_));
  AOI21_X1  g0298(.A(new_n676_), .B1(new_n467_), .B2(G124), .ZN(new_n677_));
  OR2_X1    g0299(.A1(new_n677_), .A2(G3743), .ZN(new_n678_));
  NAND2_X1  g0300(.A1(new_n677_), .A2(G3743), .ZN(new_n679_));
  NAND2_X1  g0301(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g0302(.A(new_n680_), .ZN(new_n681_));
  INV_X1    g0303(.A(G130), .ZN(new_n682_));
  NOR2_X1   g0304(.A1(new_n682_), .A2(G18), .ZN(new_n683_));
  AOI21_X1  g0305(.A(new_n683_), .B1(G18), .B2(G234), .ZN(new_n684_));
  OR2_X1    g0306(.A1(new_n684_), .A2(G3729), .ZN(new_n685_));
  NAND2_X1  g0307(.A1(new_n684_), .A2(G3729), .ZN(new_n686_));
  NAND2_X1  g0308(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g0309(.A(new_n687_), .B(KEYINPUT13), .Z(new_n688_));
  INV_X1    g0310(.A(G127), .ZN(new_n689_));
  NOR2_X1   g0311(.A1(new_n689_), .A2(G18), .ZN(new_n690_));
  AOI21_X1  g0312(.A(new_n690_), .B1(G18), .B2(G233), .ZN(new_n691_));
  NAND2_X1  g0313(.A1(new_n691_), .A2(G3737), .ZN(new_n692_));
  INV_X1    g0314(.A(new_n692_), .ZN(new_n693_));
  NOR2_X1   g0315(.A1(new_n691_), .A2(G3737), .ZN(new_n694_));
  NOR2_X1   g0316(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g0317(.A1(new_n675_), .A2(new_n681_), .A3(new_n688_), .A4(new_n695_), .ZN(new_n696_));
  INV_X1    g0318(.A(new_n678_), .ZN(new_n697_));
  XNOR2_X1  g0319(.A(new_n685_), .B(KEYINPUT14), .ZN(new_n698_));
  OAI21_X1  g0320(.A(new_n698_), .B1(G3737), .B2(new_n691_), .ZN(new_n699_));
  NAND2_X1  g0321(.A1(new_n692_), .A2(new_n679_), .ZN(new_n700_));
  INV_X1    g0322(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g0323(.A(new_n697_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g0324(.A(new_n630_), .B1(new_n696_), .B2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g0325(.A1(new_n628_), .A2(G3749), .ZN(new_n704_));
  OAI211_X1 g0326(.A(new_n590_), .B(new_n626_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g0327(.A(new_n539_), .B1(new_n547_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g0328(.A(G214), .ZN(new_n707_));
  AOI21_X1  g0329(.A(new_n454_), .B1(G18), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g0330(.A(G1480), .ZN(new_n709_));
  OR2_X1    g0331(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g0332(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g0333(.A1(new_n708_), .A2(new_n709_), .ZN(new_n712_));
  INV_X1    g0334(.A(new_n712_), .ZN(new_n713_));
  NOR2_X1   g0335(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g0336(.A(new_n714_), .ZN(new_n715_));
  INV_X1    g0337(.A(G213), .ZN(new_n716_));
  AOI21_X1  g0338(.A(new_n454_), .B1(G18), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g0339(.A(G1486), .ZN(new_n718_));
  NAND2_X1  g0340(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g0341(.A(new_n719_), .ZN(new_n720_));
  NOR2_X1   g0342(.A1(new_n717_), .A2(new_n718_), .ZN(new_n721_));
  NOR2_X1   g0343(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g0344(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g0345(.A1(new_n715_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g0346(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g0347(.A1(G1496), .A2(G4528), .ZN(new_n726_));
  XNOR2_X1  g0348(.A(new_n726_), .B(G38), .ZN(new_n727_));
  INV_X1    g0349(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g0350(.A1(G1492), .A2(G4528), .ZN(new_n729_));
  XOR2_X1   g0351(.A(new_n729_), .B(G38), .Z(new_n730_));
  NAND2_X1  g0352(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g0353(.A(G1462), .ZN(new_n732_));
  OAI211_X1 g0354(.A(new_n448_), .B(KEYINPUT4), .C1(new_n467_), .C2(G209), .ZN(new_n733_));
  INV_X1    g0355(.A(new_n733_), .ZN(new_n734_));
  INV_X1    g0356(.A(G209), .ZN(new_n735_));
  NAND2_X1  g0357(.A1(new_n735_), .A2(G18), .ZN(new_n736_));
  AOI21_X1  g0358(.A(KEYINPUT4), .B1(new_n736_), .B2(new_n448_), .ZN(new_n737_));
  OAI21_X1  g0359(.A(new_n732_), .B1(new_n734_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g0360(.A(new_n448_), .B1(new_n467_), .B2(G215), .ZN(new_n739_));
  NAND2_X1  g0361(.A1(new_n739_), .A2(G106), .ZN(new_n740_));
  INV_X1    g0362(.A(G215), .ZN(new_n741_));
  NAND2_X1  g0363(.A1(new_n741_), .A2(G18), .ZN(new_n742_));
  INV_X1    g0364(.A(G106), .ZN(new_n743_));
  NAND3_X1  g0365(.A1(new_n742_), .A2(new_n743_), .A3(new_n448_), .ZN(new_n744_));
  AND2_X1   g0366(.A1(new_n740_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g0367(.A(G1469), .ZN(new_n746_));
  OAI211_X1 g0368(.A(new_n448_), .B(new_n746_), .C1(new_n467_), .C2(G216), .ZN(new_n747_));
  INV_X1    g0369(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g0370(.A(G216), .ZN(new_n749_));
  NAND2_X1  g0371(.A1(new_n749_), .A2(G18), .ZN(new_n750_));
  AOI21_X1  g0372(.A(new_n746_), .B1(new_n750_), .B2(new_n448_), .ZN(new_n751_));
  NOR2_X1   g0373(.A1(new_n748_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g0374(.A(new_n448_), .B1(new_n467_), .B2(G209), .ZN(new_n753_));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n754_));
  NAND2_X1  g0376(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g0377(.A1(new_n755_), .A2(G1462), .A3(new_n733_), .ZN(new_n756_));
  NAND4_X1  g0378(.A1(new_n738_), .A2(new_n745_), .A3(new_n752_), .A4(new_n756_), .ZN(new_n757_));
  NOR3_X1   g0379(.A1(new_n725_), .A2(new_n731_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g0380(.A1(new_n706_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g0381(.A(new_n587_), .ZN(new_n760_));
  NOR2_X1   g0382(.A1(new_n567_), .A2(G4427), .ZN(new_n761_));
  AOI21_X1  g0383(.A(new_n761_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n762_));
  OAI21_X1  g0384(.A(new_n760_), .B1(new_n762_), .B2(new_n586_), .ZN(new_n763_));
  NAND2_X1  g0385(.A1(new_n763_), .A2(new_n581_), .ZN(new_n764_));
  INV_X1    g0386(.A(new_n578_), .ZN(new_n765_));
  AOI21_X1  g0387(.A(new_n765_), .B1(G18), .B2(G219), .ZN(new_n766_));
  OAI21_X1  g0388(.A(new_n764_), .B1(G4437), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g0389(.A(new_n609_), .ZN(new_n768_));
  NOR2_X1   g0390(.A1(new_n768_), .A2(new_n596_), .ZN(new_n769_));
  XNOR2_X1  g0391(.A(new_n769_), .B(KEYINPUT19), .ZN(new_n770_));
  INV_X1    g0392(.A(new_n616_), .ZN(new_n771_));
  NOR2_X1   g0393(.A1(new_n771_), .A2(new_n621_), .ZN(new_n772_));
  NAND3_X1  g0394(.A1(new_n604_), .A2(new_n610_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g0395(.A(G4405), .B1(new_n597_), .B2(new_n598_), .ZN(new_n774_));
  AOI21_X1  g0396(.A(new_n774_), .B1(new_n602_), .B2(new_n615_), .ZN(new_n775_));
  INV_X1    g0397(.A(new_n775_), .ZN(new_n776_));
  NAND3_X1  g0398(.A1(new_n610_), .A2(new_n595_), .A3(new_n776_), .ZN(new_n777_));
  AND4_X1   g0399(.A1(new_n594_), .A2(new_n770_), .A3(new_n773_), .A4(new_n777_), .ZN(new_n778_));
  INV_X1    g0400(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g0401(.A(new_n767_), .B1(new_n590_), .B2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g0402(.A1(new_n780_), .A2(new_n547_), .ZN(new_n781_));
  AOI22_X1  g0403(.A1(new_n781_), .A2(new_n758_), .B1(G38), .B2(new_n731_), .ZN(new_n782_));
  OAI211_X1 g0404(.A(new_n448_), .B(new_n732_), .C1(new_n467_), .C2(G209), .ZN(new_n783_));
  OR3_X1    g0405(.A1(new_n725_), .A2(KEYINPUT18), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g0406(.A(KEYINPUT18), .B1(new_n725_), .B2(new_n783_), .ZN(new_n785_));
  NAND4_X1  g0407(.A1(new_n784_), .A2(new_n745_), .A3(new_n752_), .A4(new_n785_), .ZN(new_n786_));
  NAND3_X1  g0408(.A1(new_n748_), .A2(new_n740_), .A3(new_n744_), .ZN(new_n787_));
  AOI21_X1  g0409(.A(new_n711_), .B1(new_n744_), .B2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g0410(.A1(new_n788_), .A2(new_n713_), .A3(new_n720_), .ZN(new_n789_));
  OR2_X1    g0411(.A1(new_n789_), .A2(new_n721_), .ZN(new_n790_));
  NAND2_X1  g0412(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g0413(.A(new_n791_), .ZN(new_n792_));
  OAI211_X1 g0414(.A(new_n759_), .B(new_n782_), .C1(new_n731_), .C2(new_n792_), .ZN(G246));
  NOR2_X1   g0415(.A1(G18), .A2(G110), .ZN(new_n794_));
  AOI21_X1  g0416(.A(new_n794_), .B1(G18), .B2(G2256), .ZN(new_n795_));
  INV_X1    g0417(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g0418(.A(new_n448_), .B1(new_n467_), .B2(G173), .ZN(new_n797_));
  OR2_X1    g0419(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g0420(.A1(G18), .A2(G109), .ZN(new_n799_));
  AOI21_X1  g0421(.A(new_n799_), .B1(G18), .B2(G2253), .ZN(new_n800_));
  INV_X1    g0422(.A(new_n800_), .ZN(new_n801_));
  OR2_X1    g0423(.A1(new_n467_), .A2(G174), .ZN(new_n802_));
  NAND2_X1  g0424(.A1(new_n802_), .A2(new_n448_), .ZN(new_n803_));
  AOI22_X1  g0425(.A1(new_n797_), .A2(new_n796_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g0426(.A1(G18), .A2(G86), .ZN(new_n805_));
  AOI21_X1  g0427(.A(new_n805_), .B1(G18), .B2(G2247), .ZN(new_n806_));
  INV_X1    g0428(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g0429(.A(new_n448_), .B1(new_n467_), .B2(G175), .ZN(new_n808_));
  NOR2_X1   g0430(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g0431(.A1(new_n801_), .A2(new_n803_), .ZN(new_n810_));
  OAI21_X1  g0432(.A(new_n804_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g0433(.A(new_n810_), .B1(new_n808_), .B2(new_n807_), .ZN(new_n812_));
  INV_X1    g0434(.A(new_n809_), .ZN(new_n813_));
  NAND4_X1  g0435(.A1(new_n812_), .A2(new_n804_), .A3(new_n813_), .A4(new_n798_), .ZN(new_n814_));
  OAI21_X1  g0436(.A(new_n448_), .B1(new_n467_), .B2(G176), .ZN(new_n815_));
  INV_X1    g0437(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g0438(.A1(G18), .A2(G63), .ZN(new_n817_));
  AOI21_X1  g0439(.A(new_n817_), .B1(G18), .B2(G2239), .ZN(new_n818_));
  NAND2_X1  g0440(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g0441(.A(new_n798_), .B(new_n811_), .C1(new_n814_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g0442(.A(G85), .ZN(new_n821_));
  OR3_X1    g0443(.A1(new_n821_), .A2(KEYINPUT25), .A3(G18), .ZN(new_n822_));
  OAI21_X1  g0444(.A(KEYINPUT25), .B1(new_n821_), .B2(G18), .ZN(new_n823_));
  OAI211_X1 g0445(.A(new_n822_), .B(new_n823_), .C1(new_n467_), .C2(G2230), .ZN(new_n824_));
  NAND2_X1  g0446(.A1(G18), .A2(G178), .ZN(new_n825_));
  OAI21_X1  g0447(.A(new_n825_), .B1(new_n473_), .B2(G18), .ZN(new_n826_));
  NAND2_X1  g0448(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  MUX2_X1   g0449(.A(G144), .B(G179), .S(G18), .Z(new_n828_));
  NOR2_X1   g0450(.A1(G18), .A2(G84), .ZN(new_n829_));
  AOI21_X1  g0451(.A(new_n829_), .B1(G18), .B2(G2224), .ZN(new_n830_));
  NAND2_X1  g0452(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  XOR2_X1   g0453(.A(new_n828_), .B(new_n830_), .Z(new_n832_));
  XNOR2_X1  g0454(.A(new_n832_), .B(KEYINPUT26), .ZN(new_n833_));
  INV_X1    g0455(.A(KEYINPUT27), .ZN(new_n834_));
  INV_X1    g0456(.A(G83), .ZN(new_n835_));
  OAI21_X1  g0457(.A(new_n834_), .B1(new_n835_), .B2(G18), .ZN(new_n836_));
  NAND3_X1  g0458(.A1(new_n467_), .A2(KEYINPUT27), .A3(G83), .ZN(new_n837_));
  OAI211_X1 g0459(.A(new_n836_), .B(new_n837_), .C1(new_n467_), .C2(G2218), .ZN(new_n838_));
  INV_X1    g0460(.A(G180), .ZN(new_n839_));
  OAI21_X1  g0461(.A(new_n478_), .B1(new_n467_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g0462(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g0463(.A(new_n498_), .B1(G18), .B2(G171), .ZN(new_n842_));
  NOR2_X1   g0464(.A1(G18), .A2(G65), .ZN(new_n843_));
  AOI21_X1  g0465(.A(new_n843_), .B1(G18), .B2(G2211), .ZN(new_n844_));
  INV_X1    g0466(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g0467(.A(new_n841_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g0468(.A1(new_n833_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g0469(.A1(new_n838_), .A2(new_n840_), .ZN(new_n848_));
  OAI211_X1 g0470(.A(new_n827_), .B(new_n831_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  OR2_X1    g0471(.A1(new_n824_), .A2(new_n826_), .ZN(new_n850_));
  NOR2_X1   g0472(.A1(G18), .A2(G64), .ZN(new_n851_));
  AOI21_X1  g0473(.A(new_n851_), .B1(G18), .B2(G2236), .ZN(new_n852_));
  INV_X1    g0474(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g0475(.A(new_n448_), .B1(new_n467_), .B2(G177), .ZN(new_n854_));
  NAND2_X1  g0476(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g0477(.A1(new_n849_), .A2(new_n850_), .A3(new_n855_), .ZN(new_n856_));
  OR2_X1    g0478(.A1(new_n853_), .A2(new_n854_), .ZN(new_n857_));
  NAND2_X1  g0479(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g0480(.A(new_n816_), .B(new_n818_), .ZN(new_n859_));
  NOR2_X1   g0481(.A1(new_n814_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g0482(.A(new_n820_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g0483(.A(new_n765_), .B1(G18), .B2(G189), .ZN(new_n862_));
  INV_X1    g0484(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g0485(.A1(G18), .A2(G62), .ZN(new_n864_));
  AOI21_X1  g0486(.A(new_n864_), .B1(G18), .B2(G4437), .ZN(new_n865_));
  NAND2_X1  g0487(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g0488(.A1(new_n863_), .A2(new_n865_), .ZN(new_n867_));
  AOI21_X1  g0489(.A(new_n583_), .B1(G18), .B2(G190), .ZN(new_n868_));
  INV_X1    g0490(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g0491(.A1(G18), .A2(G61), .ZN(new_n870_));
  AOI21_X1  g0492(.A(new_n870_), .B1(G18), .B2(G4432), .ZN(new_n871_));
  NAND2_X1  g0493(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g0494(.A(new_n867_), .ZN(new_n873_));
  OR2_X1    g0495(.A1(new_n869_), .A2(new_n871_), .ZN(new_n874_));
  AND4_X1   g0496(.A1(new_n873_), .A2(new_n874_), .A3(new_n872_), .A4(new_n866_), .ZN(new_n875_));
  INV_X1    g0497(.A(new_n552_), .ZN(new_n876_));
  AOI21_X1  g0498(.A(new_n876_), .B1(G18), .B2(G191), .ZN(new_n877_));
  INV_X1    g0499(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g0500(.A1(G18), .A2(G60), .ZN(new_n879_));
  AOI21_X1  g0501(.A(new_n879_), .B1(G18), .B2(G4427), .ZN(new_n880_));
  OAI21_X1  g0502(.A(new_n875_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g0503(.A(new_n572_), .B1(G18), .B2(G192), .ZN(new_n882_));
  INV_X1    g0504(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g0505(.A1(G18), .A2(G79), .ZN(new_n884_));
  AOI21_X1  g0506(.A(new_n884_), .B1(G18), .B2(G4420), .ZN(new_n885_));
  AOI22_X1  g0507(.A1(new_n878_), .A2(new_n880_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  OAI221_X1 g0508(.A(new_n866_), .B1(new_n867_), .B2(new_n872_), .C1(new_n881_), .C2(new_n886_), .ZN(new_n887_));
  INV_X1    g0509(.A(new_n611_), .ZN(new_n888_));
  AOI21_X1  g0510(.A(new_n888_), .B1(G18), .B2(G196), .ZN(new_n889_));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n890_));
  OAI21_X1  g0512(.A(new_n890_), .B1(new_n467_), .B2(G4400), .ZN(new_n891_));
  INV_X1    g0513(.A(G4400), .ZN(new_n892_));
  NAND3_X1  g0514(.A1(new_n892_), .A2(KEYINPUT30), .A3(G18), .ZN(new_n893_));
  AOI22_X1  g0515(.A1(new_n891_), .A2(new_n893_), .B1(new_n467_), .B2(G78), .ZN(new_n894_));
  NOR2_X1   g0516(.A1(new_n889_), .A2(new_n894_), .ZN(new_n895_));
  AND2_X1   g0517(.A1(new_n889_), .A2(new_n894_), .ZN(new_n896_));
  NOR2_X1   g0518(.A1(G18), .A2(G77), .ZN(new_n897_));
  AOI21_X1  g0519(.A(new_n897_), .B1(G18), .B2(G4394), .ZN(new_n898_));
  INV_X1    g0520(.A(G187), .ZN(new_n899_));
  OAI21_X1  g0521(.A(new_n617_), .B1(new_n467_), .B2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g0522(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g0523(.A1(new_n896_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g0524(.A1(G18), .A2(G59), .ZN(new_n903_));
  AOI21_X1  g0525(.A(new_n903_), .B1(G18), .B2(G4405), .ZN(new_n904_));
  XOR2_X1   g0526(.A(KEYINPUT29), .B(G195), .Z(new_n905_));
  OAI21_X1  g0527(.A(new_n597_), .B1(new_n905_), .B2(new_n467_), .ZN(new_n906_));
  AOI211_X1 g0528(.A(new_n895_), .B(new_n902_), .C1(new_n904_), .C2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g0529(.A1(new_n906_), .A2(new_n904_), .ZN(new_n908_));
  AOI21_X1  g0530(.A(new_n605_), .B1(G18), .B2(G194), .ZN(new_n909_));
  NOR2_X1   g0531(.A1(G18), .A2(G81), .ZN(new_n910_));
  AOI21_X1  g0532(.A(new_n910_), .B1(G18), .B2(G4410), .ZN(new_n911_));
  INV_X1    g0533(.A(new_n911_), .ZN(new_n912_));
  OAI22_X1  g0534(.A1(new_n907_), .A2(new_n908_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  XOR2_X1   g0535(.A(KEYINPUT28), .B(G193), .Z(new_n914_));
  OAI21_X1  g0536(.A(new_n591_), .B1(new_n914_), .B2(new_n467_), .ZN(new_n915_));
  NOR2_X1   g0537(.A1(G18), .A2(G80), .ZN(new_n916_));
  AOI21_X1  g0538(.A(new_n916_), .B1(G18), .B2(G4415), .ZN(new_n917_));
  NOR2_X1   g0539(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g0540(.A(new_n918_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n919_));
  AOI22_X1  g0541(.A1(new_n913_), .A2(new_n919_), .B1(new_n917_), .B2(new_n915_), .ZN(new_n920_));
  MUX2_X1   g0542(.A(G100), .B(G200), .S(G18), .Z(new_n921_));
  INV_X1    g0543(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g0544(.A1(G18), .A2(G3749), .ZN(new_n923_));
  OAI21_X1  g0545(.A(new_n923_), .B1(G18), .B2(G56), .ZN(new_n924_));
  OR2_X1    g0546(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g0547(.A1(G18), .A2(G202), .ZN(new_n926_));
  OAI21_X1  g0548(.A(new_n926_), .B1(new_n689_), .B2(G18), .ZN(new_n927_));
  NOR2_X1   g0549(.A1(G18), .A2(G53), .ZN(new_n928_));
  AOI21_X1  g0550(.A(new_n928_), .B1(G18), .B2(G3729), .ZN(new_n929_));
  NAND2_X1  g0551(.A1(G18), .A2(G203), .ZN(new_n930_));
  OAI21_X1  g0552(.A(new_n930_), .B1(new_n682_), .B2(G18), .ZN(new_n931_));
  AND2_X1   g0553(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g0554(.A1(G18), .A2(G3737), .ZN(new_n933_));
  OAI21_X1  g0555(.A(new_n933_), .B1(G18), .B2(G54), .ZN(new_n934_));
  INV_X1    g0556(.A(new_n934_), .ZN(new_n935_));
  OAI21_X1  g0557(.A(new_n927_), .B1(new_n932_), .B2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g0558(.A1(new_n932_), .A2(new_n935_), .ZN(new_n937_));
  MUX2_X1   g0559(.A(G124), .B(G201), .S(G18), .Z(new_n938_));
  NAND2_X1  g0560(.A1(G18), .A2(G3743), .ZN(new_n939_));
  OAI21_X1  g0561(.A(new_n939_), .B1(G18), .B2(G55), .ZN(new_n940_));
  INV_X1    g0562(.A(new_n940_), .ZN(new_n941_));
  NAND2_X1  g0563(.A1(new_n938_), .A2(new_n941_), .ZN(new_n942_));
  NAND3_X1  g0564(.A1(new_n936_), .A2(new_n937_), .A3(new_n942_), .ZN(new_n943_));
  NOR2_X1   g0565(.A1(new_n938_), .A2(new_n941_), .ZN(new_n944_));
  AOI21_X1  g0566(.A(new_n944_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n945_));
  NAND2_X1  g0567(.A1(new_n943_), .A2(new_n945_), .ZN(new_n946_));
  NAND3_X1  g0568(.A1(new_n945_), .A2(new_n925_), .A3(new_n942_), .ZN(new_n947_));
  XOR2_X1   g0569(.A(new_n934_), .B(new_n927_), .Z(new_n948_));
  NOR2_X1   g0570(.A1(new_n929_), .A2(new_n931_), .ZN(new_n949_));
  NOR4_X1   g0571(.A1(new_n947_), .A2(new_n932_), .A3(new_n948_), .A4(new_n949_), .ZN(new_n950_));
  NOR2_X1   g0572(.A1(G18), .A2(G74), .ZN(new_n951_));
  AOI21_X1  g0573(.A(new_n951_), .B1(G18), .B2(G3705), .ZN(new_n952_));
  INV_X1    g0574(.A(G207), .ZN(new_n953_));
  OAI21_X1  g0575(.A(new_n658_), .B1(new_n467_), .B2(new_n953_), .ZN(new_n954_));
  NOR2_X1   g0576(.A1(new_n952_), .A2(new_n954_), .ZN(new_n955_));
  NOR2_X1   g0577(.A1(G18), .A2(G73), .ZN(new_n956_));
  AOI21_X1  g0578(.A(new_n956_), .B1(G18), .B2(G3723), .ZN(new_n957_));
  INV_X1    g0579(.A(G204), .ZN(new_n958_));
  OAI21_X1  g0580(.A(new_n635_), .B1(new_n467_), .B2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g0581(.A1(new_n957_), .A2(new_n959_), .ZN(new_n960_));
  INV_X1    g0582(.A(G89), .ZN(new_n961_));
  NAND2_X1  g0583(.A1(new_n467_), .A2(G41), .ZN(new_n962_));
  NOR2_X1   g0584(.A1(G18), .A2(G70), .ZN(new_n963_));
  AOI21_X1  g0585(.A(new_n961_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  AOI22_X1  g0586(.A1(new_n960_), .A2(new_n964_), .B1(new_n954_), .B2(new_n952_), .ZN(new_n965_));
  NAND3_X1  g0587(.A1(new_n467_), .A2(G41), .A3(G70), .ZN(new_n966_));
  AOI21_X1  g0588(.A(new_n955_), .B1(new_n965_), .B2(new_n966_), .ZN(new_n967_));
  INV_X1    g0589(.A(G206), .ZN(new_n968_));
  OAI21_X1  g0590(.A(new_n640_), .B1(new_n467_), .B2(new_n968_), .ZN(new_n969_));
  XNOR2_X1  g0591(.A(new_n969_), .B(KEYINPUT21), .ZN(new_n970_));
  NOR2_X1   g0592(.A1(G18), .A2(G76), .ZN(new_n971_));
  AOI21_X1  g0593(.A(new_n971_), .B1(G18), .B2(G3711), .ZN(new_n972_));
  INV_X1    g0594(.A(new_n972_), .ZN(new_n973_));
  NAND2_X1  g0595(.A1(new_n970_), .A2(new_n973_), .ZN(new_n974_));
  NOR2_X1   g0596(.A1(new_n648_), .A2(G18), .ZN(new_n975_));
  AOI21_X1  g0597(.A(new_n975_), .B1(G18), .B2(G205), .ZN(new_n976_));
  INV_X1    g0598(.A(new_n976_), .ZN(new_n977_));
  INV_X1    g0599(.A(G75), .ZN(new_n978_));
  OAI21_X1  g0600(.A(KEYINPUT20), .B1(new_n978_), .B2(G18), .ZN(new_n979_));
  NOR2_X1   g0601(.A1(new_n467_), .A2(G3717), .ZN(new_n980_));
  MUX2_X1   g0602(.A(new_n979_), .B(KEYINPUT20), .S(new_n980_), .Z(new_n981_));
  AOI22_X1  g0603(.A1(new_n967_), .A2(new_n974_), .B1(new_n977_), .B2(new_n981_), .ZN(new_n982_));
  OR2_X1    g0604(.A1(new_n970_), .A2(new_n973_), .ZN(new_n983_));
  INV_X1    g0605(.A(new_n981_), .ZN(new_n984_));
  AOI22_X1  g0606(.A1(new_n982_), .A2(new_n983_), .B1(new_n976_), .B2(new_n984_), .ZN(new_n985_));
  INV_X1    g0607(.A(new_n960_), .ZN(new_n986_));
  OAI21_X1  g0608(.A(new_n950_), .B1(new_n985_), .B2(new_n986_), .ZN(new_n987_));
  NOR2_X1   g0609(.A1(new_n957_), .A2(new_n959_), .ZN(new_n988_));
  OAI211_X1 g0610(.A(new_n925_), .B(new_n946_), .C1(new_n987_), .C2(new_n988_), .ZN(new_n989_));
  NOR2_X1   g0611(.A1(new_n909_), .A2(new_n912_), .ZN(new_n990_));
  NOR4_X1   g0612(.A1(new_n908_), .A2(new_n896_), .A3(new_n895_), .A4(new_n990_), .ZN(new_n991_));
  AOI21_X1  g0613(.A(new_n918_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n992_));
  NAND3_X1  g0614(.A1(new_n989_), .A2(new_n991_), .A3(new_n992_), .ZN(new_n993_));
  NOR2_X1   g0615(.A1(new_n898_), .A2(new_n900_), .ZN(new_n994_));
  AOI21_X1  g0616(.A(new_n994_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n995_));
  NAND2_X1  g0617(.A1(new_n995_), .A2(new_n901_), .ZN(new_n996_));
  OAI21_X1  g0618(.A(new_n920_), .B1(new_n993_), .B2(new_n996_), .ZN(new_n997_));
  INV_X1    g0619(.A(new_n886_), .ZN(new_n998_));
  NOR2_X1   g0620(.A1(new_n883_), .A2(new_n885_), .ZN(new_n999_));
  NOR3_X1   g0621(.A1(new_n881_), .A2(new_n998_), .A3(new_n999_), .ZN(new_n1000_));
  AOI21_X1  g0622(.A(new_n887_), .B1(new_n997_), .B2(new_n1000_), .ZN(new_n1001_));
  INV_X1    g0623(.A(new_n842_), .ZN(new_n1002_));
  OAI21_X1  g0624(.A(new_n833_), .B1(new_n1002_), .B2(new_n844_), .ZN(new_n1003_));
  NOR3_X1   g0625(.A1(new_n1003_), .A2(new_n848_), .A3(new_n846_), .ZN(new_n1004_));
  AND3_X1   g0626(.A1(new_n857_), .A2(new_n827_), .A3(new_n855_), .ZN(new_n1005_));
  NAND4_X1  g0627(.A1(new_n1004_), .A2(new_n860_), .A3(new_n850_), .A4(new_n1005_), .ZN(new_n1006_));
  OAI21_X1  g0628(.A(new_n861_), .B1(new_n1001_), .B2(new_n1006_), .ZN(new_n1007_));
  OR2_X1    g0629(.A1(new_n467_), .A2(G169), .ZN(new_n1008_));
  NAND2_X1  g0630(.A1(new_n1008_), .A2(new_n448_), .ZN(new_n1009_));
  NAND2_X1  g0631(.A1(G18), .A2(G1469), .ZN(new_n1010_));
  OAI21_X1  g0632(.A(new_n1010_), .B1(G18), .B2(G111), .ZN(new_n1011_));
  NAND2_X1  g0633(.A1(new_n1009_), .A2(new_n1011_), .ZN(new_n1012_));
  NOR2_X1   g0634(.A1(G18), .A2(G87), .ZN(new_n1013_));
  AOI21_X1  g0635(.A(new_n1013_), .B1(G18), .B2(G106), .ZN(new_n1014_));
  OAI21_X1  g0636(.A(new_n448_), .B1(new_n467_), .B2(G168), .ZN(new_n1015_));
  XNOR2_X1  g0637(.A(new_n1014_), .B(new_n1015_), .ZN(new_n1016_));
  NOR2_X1   g0638(.A1(G18), .A2(G112), .ZN(new_n1017_));
  AOI21_X1  g0639(.A(new_n1017_), .B1(G18), .B2(G1480), .ZN(new_n1018_));
  INV_X1    g0640(.A(new_n1018_), .ZN(new_n1019_));
  OAI21_X1  g0641(.A(new_n448_), .B1(new_n467_), .B2(G167), .ZN(new_n1020_));
  NAND2_X1  g0642(.A1(new_n1019_), .A2(new_n1020_), .ZN(new_n1021_));
  AND2_X1   g0643(.A1(new_n1016_), .A2(new_n1021_), .ZN(new_n1022_));
  OR2_X1    g0644(.A1(new_n467_), .A2(G166), .ZN(new_n1023_));
  NAND2_X1  g0645(.A1(new_n1023_), .A2(new_n448_), .ZN(new_n1024_));
  NAND2_X1  g0646(.A1(G18), .A2(G1486), .ZN(new_n1025_));
  OAI21_X1  g0647(.A(new_n1025_), .B1(G18), .B2(G88), .ZN(new_n1026_));
  XNOR2_X1  g0648(.A(new_n1024_), .B(new_n1026_), .ZN(new_n1027_));
  XNOR2_X1  g0649(.A(new_n1027_), .B(KEYINPUT22), .ZN(new_n1028_));
  NOR2_X1   g0650(.A1(G18), .A2(G113), .ZN(new_n1029_));
  AOI21_X1  g0651(.A(new_n1029_), .B1(G18), .B2(G1462), .ZN(new_n1030_));
  NAND2_X1  g0652(.A1(new_n1030_), .A2(new_n448_), .ZN(new_n1031_));
  OAI21_X1  g0653(.A(new_n1031_), .B1(new_n1009_), .B2(new_n1011_), .ZN(new_n1032_));
  OR2_X1    g0654(.A1(new_n1019_), .A2(new_n1020_), .ZN(new_n1033_));
  OAI21_X1  g0655(.A(new_n1033_), .B1(new_n448_), .B2(new_n1030_), .ZN(new_n1034_));
  NOR3_X1   g0656(.A1(new_n1028_), .A2(new_n1032_), .A3(new_n1034_), .ZN(new_n1035_));
  NAND4_X1  g0657(.A1(new_n1007_), .A2(new_n1012_), .A3(new_n1022_), .A4(new_n1035_), .ZN(new_n1036_));
  NOR2_X1   g0658(.A1(new_n1024_), .A2(new_n1026_), .ZN(new_n1037_));
  NAND3_X1  g0659(.A1(new_n1016_), .A2(new_n1032_), .A3(new_n1012_), .ZN(new_n1038_));
  INV_X1    g0660(.A(new_n1014_), .ZN(new_n1039_));
  OAI211_X1 g0661(.A(new_n1038_), .B(new_n1033_), .C1(new_n1015_), .C2(new_n1039_), .ZN(new_n1040_));
  AND2_X1   g0662(.A1(new_n1040_), .A2(new_n1021_), .ZN(new_n1041_));
  INV_X1    g0663(.A(new_n1028_), .ZN(new_n1042_));
  AOI21_X1  g0664(.A(new_n1037_), .B1(new_n1041_), .B2(new_n1042_), .ZN(new_n1043_));
  NAND2_X1  g0665(.A1(new_n1036_), .A2(new_n1043_), .ZN(new_n1044_));
  INV_X1    g0666(.A(G2204), .ZN(new_n1045_));
  NAND2_X1  g0667(.A1(new_n1045_), .A2(G4528), .ZN(new_n1046_));
  XOR2_X1   g0668(.A(new_n1046_), .B(KEYINPUT24), .Z(new_n1047_));
  INV_X1    g0669(.A(new_n1047_), .ZN(new_n1048_));
  INV_X1    g0670(.A(G1455), .ZN(new_n1049_));
  NAND2_X1  g0671(.A1(new_n1049_), .A2(G4528), .ZN(new_n1050_));
  XOR2_X1   g0672(.A(new_n1050_), .B(KEYINPUT23), .Z(new_n1051_));
  NAND3_X1  g0673(.A1(new_n1048_), .A2(new_n1051_), .A3(G38), .ZN(new_n1052_));
  OR2_X1    g0674(.A1(new_n1051_), .A2(G38), .ZN(new_n1053_));
  OAI21_X1  g0675(.A(new_n1052_), .B1(new_n1053_), .B2(new_n1048_), .ZN(new_n1054_));
  NAND2_X1  g0676(.A1(new_n1044_), .A2(new_n1054_), .ZN(new_n1055_));
  OAI21_X1  g0677(.A(G38), .B1(new_n1047_), .B2(new_n1050_), .ZN(new_n1056_));
  NAND2_X1  g0678(.A1(new_n1055_), .A2(new_n1056_), .ZN(G258));
  NAND2_X1  g0679(.A1(new_n1055_), .A2(new_n1056_), .ZN(G264));
  NAND2_X1  g0680(.A1(new_n731_), .A2(G38), .ZN(new_n1059_));
  NAND2_X1  g0681(.A1(new_n705_), .A2(new_n780_), .ZN(new_n1060_));
  NAND3_X1  g0682(.A1(new_n1060_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n1061_));
  NAND2_X1  g0683(.A1(new_n1061_), .A2(new_n539_), .ZN(new_n1062_));
  NOR3_X1   g0684(.A1(new_n734_), .A2(new_n737_), .A3(new_n732_), .ZN(new_n1063_));
  AOI21_X1  g0685(.A(G1462), .B1(new_n755_), .B2(new_n733_), .ZN(new_n1064_));
  NOR2_X1   g0686(.A1(new_n1063_), .A2(new_n1064_), .ZN(new_n1065_));
  XOR2_X1   g0687(.A(new_n752_), .B(KEYINPUT31), .Z(new_n1066_));
  NAND4_X1  g0688(.A1(new_n724_), .A2(new_n745_), .A3(new_n1065_), .A4(new_n1066_), .ZN(new_n1067_));
  XOR2_X1   g0689(.A(new_n1067_), .B(KEYINPUT32), .Z(new_n1068_));
  AOI21_X1  g0690(.A(new_n791_), .B1(new_n1062_), .B2(new_n1068_), .ZN(new_n1069_));
  OAI21_X1  g0691(.A(new_n1059_), .B1(new_n1069_), .B2(new_n731_), .ZN(G270));
  NAND2_X1  g0692(.A1(new_n661_), .A2(new_n667_), .ZN(new_n1071_));
  INV_X1    g0693(.A(G3711), .ZN(new_n1072_));
  AOI21_X1  g0694(.A(new_n643_), .B1(new_n1072_), .B2(new_n642_), .ZN(new_n1073_));
  OAI211_X1 g0695(.A(new_n652_), .B(new_n1071_), .C1(new_n1073_), .C2(new_n668_), .ZN(new_n1074_));
  AND2_X1   g0696(.A1(new_n1074_), .A2(new_n651_), .ZN(new_n1075_));
  AND2_X1   g0697(.A1(new_n651_), .A2(new_n652_), .ZN(new_n1076_));
  INV_X1    g0698(.A(new_n662_), .ZN(new_n1077_));
  NAND3_X1  g0699(.A1(new_n1076_), .A2(new_n1073_), .A3(new_n1077_), .ZN(new_n1078_));
  INV_X1    g0700(.A(new_n438_), .ZN(new_n1079_));
  AOI21_X1  g0701(.A(new_n436_), .B1(new_n1079_), .B2(G4526), .ZN(new_n1080_));
  OAI21_X1  g0702(.A(new_n1075_), .B1(new_n1078_), .B2(new_n1080_), .ZN(new_n1081_));
  INV_X1    g0703(.A(new_n664_), .ZN(new_n1082_));
  XNOR2_X1  g0704(.A(new_n1081_), .B(new_n1082_), .ZN(G388));
  NAND2_X1  g0705(.A1(new_n1071_), .A2(new_n644_), .ZN(new_n1084_));
  OAI21_X1  g0706(.A(new_n1084_), .B1(new_n646_), .B2(new_n662_), .ZN(new_n1085_));
  INV_X1    g0707(.A(new_n1080_), .ZN(new_n1086_));
  INV_X1    g0708(.A(new_n1084_), .ZN(new_n1087_));
  OAI21_X1  g0709(.A(new_n1085_), .B1(new_n1086_), .B2(new_n1087_), .ZN(new_n1088_));
  XNOR2_X1  g0710(.A(new_n1088_), .B(new_n1076_), .ZN(G391));
  NOR2_X1   g0711(.A1(new_n668_), .A2(new_n643_), .ZN(new_n1090_));
  INV_X1    g0712(.A(new_n1090_), .ZN(new_n1091_));
  INV_X1    g0713(.A(new_n657_), .ZN(new_n1092_));
  OAI21_X1  g0714(.A(new_n661_), .B1(new_n1092_), .B2(new_n1080_), .ZN(new_n1093_));
  XNOR2_X1  g0715(.A(new_n1091_), .B(new_n1093_), .ZN(G394));
  XNOR2_X1  g0716(.A(new_n1086_), .B(new_n662_), .ZN(G397));
  NOR2_X1   g0717(.A1(new_n694_), .A2(new_n686_), .ZN(new_n1096_));
  OAI21_X1  g0718(.A(new_n678_), .B1(new_n1096_), .B2(new_n700_), .ZN(new_n1097_));
  NAND2_X1  g0719(.A1(new_n675_), .A2(new_n1097_), .ZN(new_n1098_));
  OAI21_X1  g0720(.A(new_n1098_), .B1(new_n702_), .B2(new_n675_), .ZN(new_n1099_));
  OR2_X1    g0721(.A1(new_n630_), .A2(new_n704_), .ZN(new_n1100_));
  XNOR2_X1  g0722(.A(new_n1099_), .B(new_n1100_), .ZN(G376));
  AND2_X1   g0723(.A1(new_n675_), .A2(new_n688_), .ZN(new_n1102_));
  OAI21_X1  g0724(.A(new_n692_), .B1(new_n1102_), .B2(new_n699_), .ZN(new_n1103_));
  XNOR2_X1  g0725(.A(new_n1103_), .B(new_n681_), .ZN(G379));
  INV_X1    g0726(.A(new_n686_), .ZN(new_n1105_));
  MUX2_X1   g0727(.A(new_n698_), .B(new_n1105_), .S(new_n675_), .Z(new_n1106_));
  XNOR2_X1  g0728(.A(new_n1106_), .B(new_n695_), .ZN(G382));
  INV_X1    g0729(.A(new_n688_), .ZN(new_n1108_));
  XNOR2_X1  g0730(.A(new_n675_), .B(new_n1108_), .ZN(G385));
  INV_X1    g0731(.A(G229), .ZN(new_n1110_));
  OAI21_X1  g0732(.A(new_n962_), .B1(new_n467_), .B2(new_n1110_), .ZN(new_n1111_));
  NAND2_X1  g0733(.A1(new_n467_), .A2(G44), .ZN(new_n1112_));
  INV_X1    g0734(.A(G239), .ZN(new_n1113_));
  OAI21_X1  g0735(.A(new_n1112_), .B1(new_n467_), .B2(new_n1113_), .ZN(new_n1114_));
  XNOR2_X1  g0736(.A(new_n1111_), .B(new_n1114_), .ZN(new_n1115_));
  XNOR2_X1  g0737(.A(new_n1115_), .B(new_n645_), .ZN(new_n1116_));
  XNOR2_X1  g0738(.A(new_n1116_), .B(new_n659_), .ZN(new_n1117_));
  NOR2_X1   g0739(.A1(new_n1117_), .A2(KEYINPUT33), .ZN(new_n1118_));
  XNOR2_X1  g0740(.A(new_n1118_), .B(new_n649_), .ZN(new_n1119_));
  XOR2_X1   g0741(.A(new_n628_), .B(new_n677_), .Z(new_n1120_));
  XNOR2_X1  g0742(.A(new_n1119_), .B(new_n1120_), .ZN(new_n1121_));
  XNOR2_X1  g0743(.A(new_n636_), .B(new_n684_), .ZN(new_n1122_));
  XNOR2_X1  g0744(.A(new_n1122_), .B(new_n691_), .ZN(new_n1123_));
  XNOR2_X1  g0745(.A(new_n1121_), .B(new_n1123_), .ZN(new_n1124_));
  XNOR2_X1  g0746(.A(new_n507_), .B(new_n480_), .ZN(new_n1125_));
  XOR2_X1   g0747(.A(new_n449_), .B(new_n475_), .Z(new_n1126_));
  XNOR2_X1  g0748(.A(new_n1125_), .B(new_n1126_), .ZN(new_n1127_));
  XNOR2_X1  g0749(.A(new_n1127_), .B(new_n490_), .ZN(new_n1128_));
  NAND3_X1  g0750(.A1(new_n456_), .A2(G18), .A3(new_n459_), .ZN(new_n1129_));
  NAND3_X1  g0751(.A1(new_n460_), .A2(G18), .A3(new_n455_), .ZN(new_n1130_));
  NAND2_X1  g0752(.A1(new_n1129_), .A2(new_n1130_), .ZN(new_n1131_));
  XNOR2_X1  g0753(.A(new_n1131_), .B(new_n469_), .ZN(new_n1132_));
  NAND2_X1  g0754(.A1(new_n467_), .A2(G141), .ZN(new_n1133_));
  INV_X1    g0755(.A(new_n1133_), .ZN(new_n1134_));
  AOI21_X1  g0756(.A(new_n1134_), .B1(G18), .B2(G161), .ZN(new_n1135_));
  XOR2_X1   g0757(.A(new_n1135_), .B(new_n499_), .Z(new_n1136_));
  XNOR2_X1  g0758(.A(new_n1132_), .B(new_n1136_), .ZN(new_n1137_));
  XNOR2_X1  g0759(.A(new_n1128_), .B(new_n1137_), .ZN(new_n1138_));
  XNOR2_X1  g0760(.A(new_n584_), .B(new_n573_), .ZN(new_n1139_));
  INV_X1    g0761(.A(new_n1139_), .ZN(new_n1140_));
  XNOR2_X1  g0762(.A(new_n606_), .B(new_n593_), .ZN(new_n1141_));
  NAND2_X1  g0763(.A1(new_n611_), .A2(new_n612_), .ZN(new_n1142_));
  XNOR2_X1  g0764(.A(new_n599_), .B(new_n1142_), .ZN(new_n1143_));
  NOR2_X1   g0765(.A1(new_n1141_), .A2(new_n1143_), .ZN(new_n1144_));
  AND2_X1   g0766(.A1(new_n1141_), .A2(new_n1143_), .ZN(new_n1145_));
  NAND2_X1  g0767(.A1(new_n467_), .A2(G115), .ZN(new_n1146_));
  INV_X1    g0768(.A(G227), .ZN(new_n1147_));
  OAI21_X1  g0769(.A(new_n1146_), .B1(new_n467_), .B2(new_n1147_), .ZN(new_n1148_));
  XNOR2_X1  g0770(.A(new_n619_), .B(new_n1148_), .ZN(new_n1149_));
  AOI21_X1  g0771(.A(new_n1144_), .B1(new_n1145_), .B2(new_n1149_), .ZN(new_n1150_));
  OAI21_X1  g0772(.A(new_n1150_), .B1(new_n1149_), .B2(new_n1145_), .ZN(new_n1151_));
  NOR2_X1   g0773(.A1(new_n1149_), .A2(KEYINPUT35), .ZN(new_n1152_));
  AOI22_X1  g0774(.A1(new_n1151_), .A2(KEYINPUT35), .B1(new_n1145_), .B2(new_n1152_), .ZN(new_n1153_));
  NOR3_X1   g0775(.A1(new_n1141_), .A2(new_n1149_), .A3(new_n1143_), .ZN(new_n1154_));
  XOR2_X1   g0776(.A(new_n1154_), .B(KEYINPUT34), .Z(new_n1155_));
  NOR2_X1   g0777(.A1(new_n1153_), .A2(new_n1155_), .ZN(new_n1156_));
  XNOR2_X1  g0778(.A(new_n558_), .B(new_n580_), .ZN(new_n1157_));
  XNOR2_X1  g0779(.A(new_n1156_), .B(new_n1157_), .ZN(new_n1158_));
  INV_X1    g0780(.A(new_n1158_), .ZN(new_n1159_));
  OAI211_X1 g0781(.A(new_n1124_), .B(new_n1138_), .C1(new_n1140_), .C2(new_n1159_), .ZN(new_n1160_));
  AOI21_X1  g0782(.A(new_n1160_), .B1(new_n1140_), .B2(new_n1159_), .ZN(new_n1161_));
  NAND3_X1  g0783(.A1(new_n708_), .A2(G18), .A3(new_n716_), .ZN(new_n1162_));
  NAND3_X1  g0784(.A1(new_n717_), .A2(G18), .A3(new_n707_), .ZN(new_n1163_));
  NAND2_X1  g0785(.A1(new_n1162_), .A2(new_n1163_), .ZN(new_n1164_));
  NAND2_X1  g0786(.A1(new_n750_), .A2(new_n448_), .ZN(new_n1165_));
  MUX2_X1   g0787(.A(new_n750_), .B(new_n1165_), .S(new_n739_), .Z(new_n1166_));
  XOR2_X1   g0788(.A(new_n1164_), .B(new_n1166_), .Z(new_n1167_));
  XNOR2_X1  g0789(.A(G211), .B(G212), .ZN(new_n1168_));
  XNOR2_X1  g0790(.A(new_n1168_), .B(new_n735_), .ZN(new_n1169_));
  NAND3_X1  g0791(.A1(new_n1169_), .A2(G18), .A3(new_n448_), .ZN(new_n1170_));
  XNOR2_X1  g0792(.A(new_n1167_), .B(new_n1170_), .ZN(new_n1171_));
  NAND2_X1  g0793(.A1(new_n1161_), .A2(new_n1171_), .ZN(G412));
  XOR2_X1   g0794(.A(new_n904_), .B(new_n898_), .Z(new_n1173_));
  XNOR2_X1  g0795(.A(new_n1173_), .B(new_n894_), .ZN(new_n1174_));
  NAND2_X1  g0796(.A1(new_n467_), .A2(G58), .ZN(new_n1175_));
  OAI21_X1  g0797(.A(new_n1175_), .B1(new_n467_), .B2(G4393), .ZN(new_n1176_));
  XNOR2_X1  g0798(.A(new_n1174_), .B(new_n1176_), .ZN(new_n1177_));
  XNOR2_X1  g0799(.A(new_n871_), .B(new_n885_), .ZN(new_n1178_));
  XNOR2_X1  g0800(.A(new_n917_), .B(new_n911_), .ZN(new_n1179_));
  XNOR2_X1  g0801(.A(new_n1178_), .B(new_n1179_), .ZN(new_n1180_));
  XNOR2_X1  g0802(.A(new_n1177_), .B(new_n1180_), .ZN(new_n1181_));
  XNOR2_X1  g0803(.A(new_n865_), .B(new_n880_), .ZN(new_n1182_));
  OR2_X1    g0804(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1183_));
  XNOR2_X1  g0805(.A(new_n1030_), .B(new_n1011_), .ZN(new_n1184_));
  NAND2_X1  g0806(.A1(G18), .A2(G1492), .ZN(new_n1185_));
  OAI21_X1  g0807(.A(new_n1185_), .B1(G18), .B2(G1455), .ZN(new_n1186_));
  XNOR2_X1  g0808(.A(new_n1014_), .B(new_n1186_), .ZN(new_n1187_));
  XNOR2_X1  g0809(.A(new_n1184_), .B(new_n1187_), .ZN(new_n1188_));
  XNOR2_X1  g0810(.A(new_n1018_), .B(new_n1026_), .ZN(new_n1189_));
  XNOR2_X1  g0811(.A(new_n1188_), .B(new_n1189_), .ZN(new_n1190_));
  NAND2_X1  g0812(.A1(new_n467_), .A2(G114), .ZN(new_n1191_));
  OAI21_X1  g0813(.A(new_n1191_), .B1(new_n467_), .B2(G1459), .ZN(new_n1192_));
  NAND2_X1  g0814(.A1(G18), .A2(G1496), .ZN(new_n1193_));
  OAI21_X1  g0815(.A(new_n1193_), .B1(G18), .B2(G2204), .ZN(new_n1194_));
  XNOR2_X1  g0816(.A(new_n1192_), .B(new_n1194_), .ZN(new_n1195_));
  XNOR2_X1  g0817(.A(new_n1190_), .B(new_n1195_), .ZN(new_n1196_));
  AOI21_X1  g0818(.A(new_n1196_), .B1(new_n1181_), .B2(new_n1182_), .ZN(new_n1197_));
  XNOR2_X1  g0819(.A(new_n924_), .B(new_n940_), .ZN(new_n1198_));
  XNOR2_X1  g0820(.A(new_n1198_), .B(new_n935_), .ZN(new_n1199_));
  AOI21_X1  g0821(.A(new_n963_), .B1(G18), .B2(G3701), .ZN(new_n1200_));
  NAND2_X1  g0822(.A1(new_n467_), .A2(G69), .ZN(new_n1201_));
  OAI21_X1  g0823(.A(new_n1201_), .B1(new_n467_), .B2(G3698), .ZN(new_n1202_));
  XNOR2_X1  g0824(.A(new_n1200_), .B(new_n1202_), .ZN(new_n1203_));
  XNOR2_X1  g0825(.A(new_n1199_), .B(new_n1203_), .ZN(new_n1204_));
  XNOR2_X1  g0826(.A(new_n1204_), .B(new_n984_), .ZN(new_n1205_));
  XNOR2_X1  g0827(.A(new_n957_), .B(new_n972_), .ZN(new_n1206_));
  XNOR2_X1  g0828(.A(new_n929_), .B(new_n952_), .ZN(new_n1207_));
  XNOR2_X1  g0829(.A(new_n1206_), .B(new_n1207_), .ZN(new_n1208_));
  XNOR2_X1  g0830(.A(new_n1205_), .B(new_n1208_), .ZN(new_n1209_));
  XNOR2_X1  g0831(.A(new_n824_), .B(new_n852_), .ZN(new_n1210_));
  NOR2_X1   g0832(.A1(new_n467_), .A2(G2208), .ZN(new_n1211_));
  AOI21_X1  g0833(.A(new_n1211_), .B1(new_n467_), .B2(G82), .ZN(new_n1212_));
  XNOR2_X1  g0834(.A(new_n1210_), .B(new_n1212_), .ZN(new_n1213_));
  XNOR2_X1  g0835(.A(new_n838_), .B(new_n800_), .ZN(new_n1214_));
  XNOR2_X1  g0836(.A(new_n1213_), .B(new_n1214_), .ZN(new_n1215_));
  XNOR2_X1  g0837(.A(new_n795_), .B(new_n806_), .ZN(new_n1216_));
  XNOR2_X1  g0838(.A(new_n1216_), .B(new_n818_), .ZN(new_n1217_));
  XNOR2_X1  g0839(.A(new_n830_), .B(new_n844_), .ZN(new_n1218_));
  XNOR2_X1  g0840(.A(new_n1217_), .B(new_n1218_), .ZN(new_n1219_));
  XNOR2_X1  g0841(.A(new_n1215_), .B(new_n1219_), .ZN(new_n1220_));
  NAND4_X1  g0842(.A1(new_n1183_), .A2(new_n1197_), .A3(new_n1209_), .A4(new_n1220_), .ZN(G414));
  XNOR2_X1  g0843(.A(new_n970_), .B(new_n976_), .ZN(new_n1222_));
  XNOR2_X1  g0844(.A(new_n1222_), .B(new_n954_), .ZN(new_n1223_));
  INV_X1    g0845(.A(new_n1112_), .ZN(new_n1224_));
  AOI21_X1  g0846(.A(new_n1224_), .B1(G18), .B2(G208), .ZN(new_n1225_));
  XNOR2_X1  g0847(.A(new_n1223_), .B(new_n1225_), .ZN(new_n1226_));
  XNOR2_X1  g0848(.A(new_n938_), .B(new_n931_), .ZN(new_n1227_));
  XNOR2_X1  g0849(.A(new_n1226_), .B(new_n1227_), .ZN(new_n1228_));
  INV_X1    g0850(.A(G198), .ZN(new_n1229_));
  OAI21_X1  g0851(.A(new_n962_), .B1(new_n467_), .B2(new_n1229_), .ZN(new_n1230_));
  XNOR2_X1  g0852(.A(new_n959_), .B(new_n1230_), .ZN(new_n1231_));
  XNOR2_X1  g0853(.A(new_n921_), .B(new_n927_), .ZN(new_n1232_));
  XNOR2_X1  g0854(.A(new_n1231_), .B(new_n1232_), .ZN(new_n1233_));
  XNOR2_X1  g0855(.A(new_n1228_), .B(new_n1233_), .ZN(new_n1234_));
  INV_X1    g0856(.A(new_n808_), .ZN(new_n1235_));
  OAI21_X1  g0857(.A(new_n1235_), .B1(new_n467_), .B2(G176), .ZN(new_n1236_));
  OAI21_X1  g0858(.A(new_n1236_), .B1(new_n816_), .B2(new_n1235_), .ZN(new_n1237_));
  XNOR2_X1  g0859(.A(new_n1237_), .B(new_n826_), .ZN(new_n1238_));
  XOR2_X1   g0860(.A(new_n828_), .B(new_n854_), .Z(new_n1239_));
  XNOR2_X1  g0861(.A(new_n1238_), .B(new_n1239_), .ZN(new_n1240_));
  MUX2_X1   g0862(.A(new_n802_), .B(new_n803_), .S(new_n797_), .Z(new_n1241_));
  XOR2_X1   g0863(.A(KEYINPUT36), .B(G181), .Z(new_n1242_));
  AOI21_X1  g0864(.A(new_n1134_), .B1(new_n1242_), .B2(G18), .ZN(new_n1243_));
  XNOR2_X1  g0865(.A(new_n1241_), .B(new_n1243_), .ZN(new_n1244_));
  XNOR2_X1  g0866(.A(new_n1240_), .B(new_n1244_), .ZN(new_n1245_));
  XOR2_X1   g0867(.A(new_n842_), .B(new_n840_), .Z(new_n1246_));
  XNOR2_X1  g0868(.A(new_n1245_), .B(new_n1246_), .ZN(new_n1247_));
  XNOR2_X1  g0869(.A(new_n862_), .B(new_n877_), .ZN(new_n1248_));
  XNOR2_X1  g0870(.A(new_n1248_), .B(new_n882_), .ZN(new_n1249_));
  XNOR2_X1  g0871(.A(new_n889_), .B(new_n909_), .ZN(new_n1250_));
  XNOR2_X1  g0872(.A(new_n1249_), .B(new_n1250_), .ZN(new_n1251_));
  INV_X1    g0873(.A(G197), .ZN(new_n1252_));
  OAI21_X1  g0874(.A(new_n1146_), .B1(new_n467_), .B2(new_n1252_), .ZN(new_n1253_));
  XOR2_X1   g0875(.A(new_n900_), .B(new_n1253_), .Z(new_n1254_));
  XNOR2_X1  g0876(.A(new_n1254_), .B(new_n915_), .ZN(new_n1255_));
  XNOR2_X1  g0877(.A(new_n906_), .B(new_n868_), .ZN(new_n1256_));
  XNOR2_X1  g0878(.A(new_n1255_), .B(new_n1256_), .ZN(new_n1257_));
  XNOR2_X1  g0879(.A(new_n1251_), .B(new_n1257_), .ZN(new_n1258_));
  MUX2_X1   g0880(.A(new_n1008_), .B(new_n1009_), .S(new_n1015_), .Z(new_n1259_));
  INV_X1    g0881(.A(new_n1259_), .ZN(new_n1260_));
  MUX2_X1   g0882(.A(new_n1023_), .B(new_n1024_), .S(new_n1020_), .Z(new_n1261_));
  OR2_X1    g0883(.A1(new_n1260_), .A2(new_n1261_), .ZN(new_n1262_));
  NAND2_X1  g0884(.A1(new_n1260_), .A2(new_n1261_), .ZN(new_n1263_));
  NAND3_X1  g0885(.A1(new_n1262_), .A2(new_n1263_), .A3(KEYINPUT37), .ZN(new_n1264_));
  XOR2_X1   g0886(.A(G164), .B(G165), .Z(new_n1265_));
  NAND3_X1  g0887(.A1(new_n1265_), .A2(G18), .A3(new_n448_), .ZN(new_n1266_));
  NOR3_X1   g0888(.A1(new_n454_), .A2(new_n467_), .A3(G170), .ZN(new_n1267_));
  XNOR2_X1  g0889(.A(new_n1266_), .B(new_n1267_), .ZN(new_n1268_));
  XNOR2_X1  g0890(.A(new_n1264_), .B(new_n1268_), .ZN(new_n1269_));
  NAND4_X1  g0891(.A1(new_n1234_), .A2(new_n1247_), .A3(new_n1258_), .A4(new_n1269_), .ZN(G416));
  NAND2_X1  g0892(.A1(G258), .A2(KEYINPUT38), .ZN(new_n1271_));
  INV_X1    g0893(.A(KEYINPUT38), .ZN(new_n1272_));
  NAND3_X1  g0894(.A1(new_n1055_), .A2(new_n1272_), .A3(new_n1056_), .ZN(new_n1273_));
  NAND2_X1  g0895(.A1(new_n1271_), .A2(new_n1273_), .ZN(G249));
  XNOR2_X1  g0896(.A(new_n1060_), .B(new_n541_), .ZN(G295));
  OR2_X1    g0897(.A1(new_n706_), .A2(new_n781_), .ZN(new_n1276_));
  INV_X1    g0898(.A(new_n1065_), .ZN(new_n1277_));
  XNOR2_X1  g0899(.A(new_n1276_), .B(new_n1277_), .ZN(G324));
  XOR2_X1   g0900(.A(new_n1001_), .B(KEYINPUT39), .Z(G252));
  OAI21_X1  g0901(.A(new_n1059_), .B1(new_n1069_), .B2(new_n731_), .ZN(G276));
  INV_X1    g0902(.A(KEYINPUT40), .ZN(new_n1281_));
  XNOR2_X1  g0903(.A(new_n514_), .B(new_n1281_), .ZN(new_n1282_));
  NAND2_X1  g0904(.A1(new_n505_), .A2(new_n1282_), .ZN(new_n1283_));
  NAND2_X1  g0905(.A1(new_n1060_), .A2(new_n542_), .ZN(new_n1284_));
  NOR2_X1   g0906(.A1(new_n1284_), .A2(new_n510_), .ZN(new_n1285_));
  AOI21_X1  g0907(.A(G2224), .B1(new_n488_), .B2(new_n489_), .ZN(new_n1286_));
  AOI21_X1  g0908(.A(new_n493_), .B1(new_n467_), .B2(G144), .ZN(new_n1287_));
  NOR2_X1   g0909(.A1(new_n1286_), .A2(new_n1287_), .ZN(new_n1288_));
  AOI21_X1  g0910(.A(new_n1283_), .B1(new_n1285_), .B2(new_n1288_), .ZN(new_n1289_));
  INV_X1    g0911(.A(new_n544_), .ZN(new_n1290_));
  XNOR2_X1  g0912(.A(new_n1289_), .B(new_n1290_), .ZN(G310));
  INV_X1    g0913(.A(new_n1287_), .ZN(new_n1292_));
  AOI21_X1  g0914(.A(new_n1286_), .B1(new_n513_), .B2(new_n1292_), .ZN(new_n1293_));
  INV_X1    g0915(.A(new_n495_), .ZN(new_n1294_));
  OAI211_X1 g0916(.A(new_n502_), .B(new_n1293_), .C1(new_n1284_), .C2(new_n1294_), .ZN(new_n1295_));
  XNOR2_X1  g0917(.A(new_n1295_), .B(new_n510_), .ZN(G313));
  NAND2_X1  g0918(.A1(new_n480_), .A2(G2218), .ZN(new_n1297_));
  INV_X1    g0919(.A(new_n1297_), .ZN(new_n1298_));
  AOI21_X1  g0920(.A(new_n1298_), .B1(new_n500_), .B2(new_n512_), .ZN(new_n1299_));
  INV_X1    g0921(.A(new_n1299_), .ZN(new_n1300_));
  NAND2_X1  g0922(.A1(new_n1284_), .A2(new_n1300_), .ZN(new_n1301_));
  INV_X1    g0923(.A(new_n1288_), .ZN(new_n1302_));
  XNOR2_X1  g0924(.A(new_n1301_), .B(new_n1302_), .ZN(G316));
  AND2_X1   g0925(.A1(new_n705_), .A2(new_n780_), .ZN(new_n1304_));
  OAI21_X1  g0926(.A(new_n500_), .B1(new_n1304_), .B2(new_n541_), .ZN(new_n1305_));
  XNOR2_X1  g0927(.A(new_n1305_), .B(new_n486_), .ZN(G319));
  INV_X1    g0928(.A(new_n751_), .ZN(new_n1307_));
  INV_X1    g0929(.A(new_n783_), .ZN(new_n1308_));
  OAI21_X1  g0930(.A(new_n1307_), .B1(new_n748_), .B2(new_n1308_), .ZN(new_n1309_));
  INV_X1    g0931(.A(new_n740_), .ZN(new_n1310_));
  OAI211_X1 g0932(.A(new_n712_), .B(new_n744_), .C1(new_n1309_), .C2(new_n1310_), .ZN(new_n1311_));
  NAND2_X1  g0933(.A1(new_n1311_), .A2(new_n710_), .ZN(new_n1312_));
  NAND3_X1  g0934(.A1(new_n1276_), .A2(new_n745_), .A3(new_n1065_), .ZN(new_n1313_));
  NAND2_X1  g0935(.A1(new_n1066_), .A2(new_n714_), .ZN(new_n1314_));
  OAI21_X1  g0936(.A(new_n1312_), .B1(new_n1313_), .B2(new_n1314_), .ZN(new_n1315_));
  XNOR2_X1  g0937(.A(new_n1315_), .B(new_n723_), .ZN(G327));
  NAND2_X1  g0938(.A1(new_n787_), .A2(KEYINPUT41), .ZN(new_n1317_));
  INV_X1    g0939(.A(KEYINPUT41), .ZN(new_n1318_));
  NAND4_X1  g0940(.A1(new_n748_), .A2(new_n740_), .A3(new_n1318_), .A4(new_n744_), .ZN(new_n1319_));
  NAND3_X1  g0941(.A1(new_n1317_), .A2(new_n744_), .A3(new_n1319_), .ZN(new_n1320_));
  INV_X1    g0942(.A(new_n1320_), .ZN(new_n1321_));
  AOI21_X1  g0943(.A(new_n1308_), .B1(new_n1276_), .B2(new_n1065_), .ZN(new_n1322_));
  NAND4_X1  g0944(.A1(new_n1307_), .A2(new_n740_), .A3(new_n744_), .A4(new_n747_), .ZN(new_n1323_));
  OAI21_X1  g0945(.A(new_n1321_), .B1(new_n1322_), .B2(new_n1323_), .ZN(new_n1324_));
  XNOR2_X1  g0946(.A(new_n1324_), .B(new_n715_), .ZN(G330));
  NAND3_X1  g0947(.A1(new_n1276_), .A2(new_n1307_), .A3(new_n1065_), .ZN(new_n1326_));
  NAND2_X1  g0948(.A1(new_n1326_), .A2(new_n1309_), .ZN(new_n1327_));
  INV_X1    g0949(.A(new_n745_), .ZN(new_n1328_));
  XNOR2_X1  g0950(.A(new_n1327_), .B(new_n1328_), .ZN(G333));
  XNOR2_X1  g0951(.A(new_n1322_), .B(new_n752_), .ZN(G336));
  NOR2_X1   g0952(.A1(G416), .A2(G414), .ZN(new_n1331_));
  NOR4_X1   g0953(.A1(G404), .A2(G406), .A3(G408), .A4(G410), .ZN(new_n1332_));
  NAND4_X1  g0954(.A1(new_n1161_), .A2(new_n1171_), .A3(new_n1331_), .A4(new_n1332_), .ZN(G418));
  OAI211_X1 g0955(.A(new_n759_), .B(new_n782_), .C1(new_n731_), .C2(new_n792_), .ZN(G273));
  AND2_X1   g0956(.A1(new_n1060_), .A2(new_n546_), .ZN(new_n1335_));
  NOR2_X1   g0957(.A1(new_n1335_), .A2(new_n517_), .ZN(new_n1336_));
  INV_X1    g0958(.A(new_n1336_), .ZN(new_n1337_));
  NAND2_X1  g0959(.A1(new_n1337_), .A2(new_n534_), .ZN(new_n1338_));
  OAI21_X1  g0960(.A(new_n1338_), .B1(new_n466_), .B2(new_n1337_), .ZN(new_n1339_));
  XNOR2_X1  g0961(.A(new_n1339_), .B(new_n535_), .ZN(G298));
  INV_X1    g0962(.A(new_n465_), .ZN(new_n1341_));
  NAND2_X1  g0963(.A1(new_n453_), .A2(new_n464_), .ZN(new_n1342_));
  NAND3_X1  g0964(.A1(new_n1336_), .A2(new_n1341_), .A3(new_n1342_), .ZN(new_n1343_));
  XOR2_X1   g0965(.A(new_n1343_), .B(KEYINPUT42), .Z(new_n1344_));
  OAI211_X1 g0966(.A(new_n1337_), .B(new_n533_), .C1(new_n532_), .C2(new_n1342_), .ZN(new_n1345_));
  NAND2_X1  g0967(.A1(new_n1344_), .A2(new_n1345_), .ZN(G301));
  OAI21_X1  g0968(.A(new_n458_), .B1(new_n1336_), .B2(new_n518_), .ZN(new_n1347_));
  XOR2_X1   g0969(.A(new_n1347_), .B(new_n526_), .Z(G304));
  XNOR2_X1  g0970(.A(new_n1336_), .B(new_n528_), .ZN(G307));
  NOR2_X1   g0971(.A1(new_n703_), .A2(new_n704_), .ZN(new_n1350_));
  XNOR2_X1  g0972(.A(new_n1350_), .B(new_n624_), .ZN(G344));
  NOR2_X1   g0973(.A1(new_n725_), .A2(new_n757_), .ZN(new_n1352_));
  AOI21_X1  g0974(.A(new_n791_), .B1(new_n1276_), .B2(new_n1352_), .ZN(new_n1353_));
  AOI21_X1  g0975(.A(G38), .B1(G1492), .B2(G4528), .ZN(new_n1354_));
  XOR2_X1   g0976(.A(new_n1354_), .B(new_n726_), .Z(new_n1355_));
  NOR2_X1   g0977(.A1(new_n1353_), .A2(new_n1355_), .ZN(new_n1356_));
  NAND2_X1  g0978(.A1(new_n729_), .A2(G38), .ZN(new_n1357_));
  XNOR2_X1  g0979(.A(new_n727_), .B(new_n1357_), .ZN(new_n1358_));
  INV_X1    g0980(.A(new_n1358_), .ZN(new_n1359_));
  AOI211_X1 g0981(.A(new_n791_), .B(new_n1359_), .C1(new_n1276_), .C2(new_n1352_), .ZN(new_n1360_));
  NOR2_X1   g0982(.A1(new_n1356_), .A2(new_n1360_), .ZN(G422));
  INV_X1    g0983(.A(KEYINPUT43), .ZN(new_n1362_));
  OAI21_X1  g0984(.A(new_n1362_), .B1(new_n1356_), .B2(new_n1360_), .ZN(new_n1363_));
  NAND2_X1  g0985(.A1(new_n1353_), .A2(new_n1358_), .ZN(new_n1364_));
  OAI211_X1 g0986(.A(new_n1364_), .B(KEYINPUT43), .C1(new_n1353_), .C2(new_n1355_), .ZN(new_n1365_));
  NAND2_X1  g0987(.A1(new_n1363_), .A2(new_n1365_), .ZN(G469));
  XNOR2_X1  g0988(.A(new_n1353_), .B(new_n730_), .ZN(G419));
  XNOR2_X1  g0989(.A(new_n1353_), .B(new_n730_), .ZN(G471));
  INV_X1    g0990(.A(new_n1350_), .ZN(new_n1369_));
  NAND4_X1  g0991(.A1(new_n1369_), .A2(new_n602_), .A3(new_n616_), .A4(new_n624_), .ZN(new_n1370_));
  NAND2_X1  g0992(.A1(new_n624_), .A2(new_n775_), .ZN(new_n1371_));
  NAND2_X1  g0993(.A1(new_n1142_), .A2(new_n892_), .ZN(new_n1372_));
  NAND3_X1  g0994(.A1(new_n1372_), .A2(new_n613_), .A3(new_n622_), .ZN(new_n1373_));
  OAI21_X1  g0995(.A(new_n775_), .B1(new_n1373_), .B2(new_n603_), .ZN(new_n1374_));
  NAND2_X1  g0996(.A1(new_n1371_), .A2(new_n1374_), .ZN(new_n1375_));
  NAND2_X1  g0997(.A1(new_n1370_), .A2(new_n1375_), .ZN(new_n1376_));
  AOI21_X1  g0998(.A(new_n609_), .B1(new_n1376_), .B2(new_n607_), .ZN(new_n1377_));
  INV_X1    g0999(.A(new_n596_), .ZN(new_n1378_));
  XNOR2_X1  g1000(.A(new_n1377_), .B(new_n1378_), .ZN(G359));
  INV_X1    g1001(.A(new_n610_), .ZN(new_n1380_));
  XNOR2_X1  g1002(.A(new_n1376_), .B(new_n1380_), .ZN(G362));
  INV_X1    g1003(.A(new_n622_), .ZN(new_n1382_));
  OAI21_X1  g1004(.A(new_n621_), .B1(new_n1350_), .B2(new_n1382_), .ZN(new_n1383_));
  AOI21_X1  g1005(.A(new_n615_), .B1(new_n1383_), .B2(new_n613_), .ZN(new_n1384_));
  INV_X1    g1006(.A(new_n603_), .ZN(new_n1385_));
  XNOR2_X1  g1007(.A(new_n1384_), .B(new_n1385_), .ZN(G365));
  XNOR2_X1  g1008(.A(new_n1383_), .B(new_n771_), .ZN(G368));
  NAND2_X1  g1009(.A1(new_n1369_), .A2(new_n626_), .ZN(new_n1388_));
  NAND2_X1  g1010(.A1(new_n1388_), .A2(new_n778_), .ZN(new_n1389_));
  INV_X1    g1011(.A(new_n581_), .ZN(new_n1390_));
  XNOR2_X1  g1012(.A(new_n763_), .B(new_n1390_), .ZN(new_n1391_));
  AOI21_X1  g1013(.A(new_n1389_), .B1(KEYINPUT44), .B2(new_n1391_), .ZN(new_n1392_));
  OAI21_X1  g1014(.A(new_n1392_), .B1(KEYINPUT44), .B2(new_n1391_), .ZN(new_n1393_));
  INV_X1    g1015(.A(new_n1389_), .ZN(new_n1394_));
  AOI21_X1  g1016(.A(new_n575_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n1395_));
  OAI21_X1  g1017(.A(new_n585_), .B1(new_n1395_), .B2(new_n761_), .ZN(new_n1396_));
  NAND2_X1  g1018(.A1(new_n1396_), .A2(new_n760_), .ZN(new_n1397_));
  XNOR2_X1  g1019(.A(new_n1397_), .B(new_n581_), .ZN(new_n1398_));
  OAI21_X1  g1020(.A(new_n1393_), .B1(new_n1394_), .B2(new_n1398_), .ZN(G347));
  OAI21_X1  g1021(.A(new_n1389_), .B1(new_n761_), .B2(new_n1395_), .ZN(new_n1400_));
  OAI21_X1  g1022(.A(new_n1400_), .B1(new_n762_), .B2(new_n1389_), .ZN(new_n1401_));
  INV_X1    g1023(.A(new_n588_), .ZN(new_n1402_));
  XNOR2_X1  g1024(.A(new_n1401_), .B(new_n1402_), .ZN(G350));
  AOI21_X1  g1025(.A(new_n576_), .B1(new_n1389_), .B2(new_n574_), .ZN(new_n1404_));
  XNOR2_X1  g1026(.A(new_n1404_), .B(new_n571_), .ZN(G353));
  INV_X1    g1027(.A(new_n577_), .ZN(new_n1406_));
  XNOR2_X1  g1028(.A(new_n1389_), .B(new_n1406_), .ZN(G356));
  INV_X1    g1029(.A(new_n496_), .ZN(new_n1408_));
  NAND2_X1  g1030(.A1(new_n497_), .A2(new_n540_), .ZN(new_n1409_));
  NAND2_X1  g1031(.A1(new_n1409_), .A2(new_n1293_), .ZN(new_n1410_));
  XNOR2_X1  g1032(.A(new_n1410_), .B(new_n544_), .ZN(new_n1411_));
  XNOR2_X1  g1033(.A(new_n486_), .B(new_n500_), .ZN(new_n1412_));
  NAND2_X1  g1034(.A1(new_n540_), .A2(KEYINPUT46), .ZN(new_n1413_));
  XNOR2_X1  g1035(.A(new_n1412_), .B(new_n1413_), .ZN(new_n1414_));
  INV_X1    g1036(.A(new_n1414_), .ZN(new_n1415_));
  NAND3_X1  g1037(.A1(new_n505_), .A2(new_n1282_), .A3(new_n543_), .ZN(new_n1416_));
  OAI21_X1  g1038(.A(new_n1300_), .B1(new_n486_), .B2(new_n541_), .ZN(new_n1417_));
  XNOR2_X1  g1039(.A(new_n1417_), .B(KEYINPUT47), .ZN(new_n1418_));
  INV_X1    g1040(.A(new_n1418_), .ZN(new_n1419_));
  NAND2_X1  g1041(.A1(new_n1416_), .A2(new_n1419_), .ZN(new_n1420_));
  NAND4_X1  g1042(.A1(new_n505_), .A2(new_n1282_), .A3(new_n1418_), .A4(new_n543_), .ZN(new_n1421_));
  AOI21_X1  g1043(.A(new_n1415_), .B1(new_n1420_), .B2(new_n1421_), .ZN(new_n1422_));
  INV_X1    g1044(.A(new_n1422_), .ZN(new_n1423_));
  NAND3_X1  g1045(.A1(new_n1420_), .A2(new_n1415_), .A3(new_n1421_), .ZN(new_n1424_));
  AOI21_X1  g1046(.A(new_n1411_), .B1(new_n1423_), .B2(new_n1424_), .ZN(new_n1425_));
  INV_X1    g1047(.A(new_n1424_), .ZN(new_n1426_));
  INV_X1    g1048(.A(new_n1411_), .ZN(new_n1427_));
  NOR3_X1   g1049(.A1(new_n1426_), .A2(new_n1427_), .A3(new_n1422_), .ZN(new_n1428_));
  OAI21_X1  g1050(.A(new_n1408_), .B1(new_n1425_), .B2(new_n1428_), .ZN(new_n1429_));
  INV_X1    g1051(.A(new_n510_), .ZN(new_n1430_));
  OAI21_X1  g1052(.A(new_n1427_), .B1(new_n1426_), .B2(new_n1422_), .ZN(new_n1431_));
  NAND3_X1  g1053(.A1(new_n1423_), .A2(new_n1411_), .A3(new_n1424_), .ZN(new_n1432_));
  NAND3_X1  g1054(.A1(new_n1431_), .A2(new_n1432_), .A3(new_n1302_), .ZN(new_n1433_));
  AND3_X1   g1055(.A1(new_n1429_), .A2(new_n1430_), .A3(new_n1433_), .ZN(new_n1434_));
  AOI21_X1  g1056(.A(new_n1430_), .B1(new_n1429_), .B2(new_n1433_), .ZN(new_n1435_));
  OAI21_X1  g1057(.A(new_n1060_), .B1(new_n1434_), .B2(new_n1435_), .ZN(new_n1436_));
  NAND2_X1  g1058(.A1(new_n1299_), .A2(new_n1292_), .ZN(new_n1437_));
  AOI21_X1  g1059(.A(new_n500_), .B1(new_n1437_), .B2(new_n492_), .ZN(new_n1438_));
  AND2_X1   g1060(.A1(new_n1293_), .A2(new_n500_), .ZN(new_n1439_));
  NOR2_X1   g1061(.A1(new_n1438_), .A2(new_n1439_), .ZN(new_n1440_));
  XOR2_X1   g1062(.A(new_n486_), .B(new_n541_), .Z(new_n1441_));
  XNOR2_X1  g1063(.A(new_n1440_), .B(new_n1441_), .ZN(new_n1442_));
  NAND2_X1  g1064(.A1(new_n1442_), .A2(new_n1300_), .ZN(new_n1443_));
  INV_X1    g1065(.A(new_n1443_), .ZN(new_n1444_));
  NOR2_X1   g1066(.A1(new_n1442_), .A2(new_n1300_), .ZN(new_n1445_));
  NAND2_X1  g1067(.A1(new_n1283_), .A2(new_n1290_), .ZN(new_n1446_));
  INV_X1    g1068(.A(new_n1446_), .ZN(new_n1447_));
  NAND3_X1  g1069(.A1(new_n505_), .A2(new_n1282_), .A3(new_n544_), .ZN(new_n1448_));
  INV_X1    g1070(.A(new_n1448_), .ZN(new_n1449_));
  OAI22_X1  g1071(.A1(new_n1444_), .A2(new_n1445_), .B1(new_n1447_), .B2(new_n1449_), .ZN(new_n1450_));
  OR2_X1    g1072(.A1(new_n1442_), .A2(new_n1300_), .ZN(new_n1451_));
  NAND4_X1  g1073(.A1(new_n1451_), .A2(new_n1446_), .A3(new_n1448_), .A4(new_n1443_), .ZN(new_n1452_));
  NAND3_X1  g1074(.A1(new_n1450_), .A2(new_n1452_), .A3(new_n496_), .ZN(new_n1453_));
  INV_X1    g1075(.A(new_n1453_), .ZN(new_n1454_));
  AOI21_X1  g1076(.A(new_n1302_), .B1(new_n1450_), .B2(new_n1452_), .ZN(new_n1455_));
  OAI211_X1 g1077(.A(KEYINPUT48), .B(new_n510_), .C1(new_n1454_), .C2(new_n1455_), .ZN(new_n1456_));
  INV_X1    g1078(.A(new_n1455_), .ZN(new_n1457_));
  OR2_X1    g1079(.A1(new_n510_), .A2(KEYINPUT48), .ZN(new_n1458_));
  NAND2_X1  g1080(.A1(new_n510_), .A2(KEYINPUT48), .ZN(new_n1459_));
  NAND4_X1  g1081(.A1(new_n1457_), .A2(new_n1453_), .A3(new_n1458_), .A4(new_n1459_), .ZN(new_n1460_));
  NAND2_X1  g1082(.A1(new_n1456_), .A2(new_n1460_), .ZN(new_n1461_));
  NAND2_X1  g1083(.A1(new_n1060_), .A2(KEYINPUT45), .ZN(new_n1462_));
  INV_X1    g1084(.A(KEYINPUT45), .ZN(new_n1463_));
  NAND2_X1  g1085(.A1(new_n1304_), .A2(new_n1463_), .ZN(new_n1464_));
  NAND3_X1  g1086(.A1(new_n1461_), .A2(new_n1462_), .A3(new_n1464_), .ZN(new_n1465_));
  NAND2_X1  g1087(.A1(new_n1436_), .A2(new_n1465_), .ZN(new_n1466_));
  NAND2_X1  g1088(.A1(new_n1464_), .A2(new_n1462_), .ZN(new_n1467_));
  NAND2_X1  g1089(.A1(new_n1467_), .A2(new_n545_), .ZN(new_n1468_));
  NAND2_X1  g1090(.A1(new_n1341_), .A2(new_n452_), .ZN(new_n1469_));
  OAI21_X1  g1091(.A(new_n463_), .B1(new_n458_), .B2(new_n520_), .ZN(new_n1470_));
  XNOR2_X1  g1092(.A(new_n1469_), .B(new_n1470_), .ZN(new_n1471_));
  XOR2_X1   g1093(.A(new_n1471_), .B(new_n535_), .Z(new_n1472_));
  AOI21_X1  g1094(.A(new_n517_), .B1(new_n1472_), .B2(new_n530_), .ZN(new_n1473_));
  OR2_X1    g1095(.A1(new_n1472_), .A2(new_n530_), .ZN(new_n1474_));
  NAND4_X1  g1096(.A1(new_n1468_), .A2(new_n1464_), .A3(new_n1473_), .A4(new_n1474_), .ZN(new_n1475_));
  XOR2_X1   g1097(.A(new_n531_), .B(new_n536_), .Z(new_n1476_));
  INV_X1    g1098(.A(new_n545_), .ZN(new_n1477_));
  NOR2_X1   g1099(.A1(new_n1304_), .A2(new_n1477_), .ZN(new_n1478_));
  OAI211_X1 g1100(.A(new_n1464_), .B(new_n1476_), .C1(new_n1478_), .C2(new_n517_), .ZN(new_n1479_));
  AND2_X1   g1101(.A1(new_n1475_), .A2(new_n1479_), .ZN(new_n1480_));
  AOI22_X1  g1102(.A1(new_n1475_), .A2(new_n1479_), .B1(new_n1461_), .B2(new_n1304_), .ZN(new_n1481_));
  NOR3_X1   g1103(.A1(new_n1425_), .A2(new_n1428_), .A3(new_n496_), .ZN(new_n1482_));
  AOI21_X1  g1104(.A(new_n1288_), .B1(new_n1431_), .B2(new_n1432_), .ZN(new_n1483_));
  NOR3_X1   g1105(.A1(new_n1482_), .A2(new_n1430_), .A3(new_n1483_), .ZN(new_n1484_));
  OAI21_X1  g1106(.A(new_n1467_), .B1(new_n1484_), .B2(new_n1434_), .ZN(new_n1485_));
  AOI22_X1  g1107(.A1(new_n1466_), .A2(new_n1480_), .B1(new_n1481_), .B2(new_n1485_), .ZN(G321));
  INV_X1    g1108(.A(new_n1066_), .ZN(new_n1487_));
  AOI21_X1  g1109(.A(new_n751_), .B1(new_n747_), .B2(new_n783_), .ZN(new_n1488_));
  NAND4_X1  g1110(.A1(new_n1317_), .A2(new_n744_), .A3(new_n1323_), .A4(new_n1319_), .ZN(new_n1489_));
  NAND2_X1  g1111(.A1(new_n1489_), .A2(new_n1308_), .ZN(new_n1490_));
  NAND4_X1  g1112(.A1(new_n1317_), .A2(new_n744_), .A3(new_n783_), .A4(new_n1319_), .ZN(new_n1491_));
  AND3_X1   g1113(.A1(new_n1490_), .A2(new_n1277_), .A3(new_n1491_), .ZN(new_n1492_));
  AOI21_X1  g1114(.A(new_n1277_), .B1(new_n1490_), .B2(new_n1491_), .ZN(new_n1493_));
  OAI21_X1  g1115(.A(new_n1488_), .B1(new_n1492_), .B2(new_n1493_), .ZN(new_n1494_));
  NAND2_X1  g1116(.A1(new_n1490_), .A2(new_n1491_), .ZN(new_n1495_));
  NAND2_X1  g1117(.A1(new_n1495_), .A2(new_n1065_), .ZN(new_n1496_));
  NAND3_X1  g1118(.A1(new_n1490_), .A2(new_n1277_), .A3(new_n1491_), .ZN(new_n1497_));
  NAND3_X1  g1119(.A1(new_n1496_), .A2(new_n1309_), .A3(new_n1497_), .ZN(new_n1498_));
  INV_X1    g1120(.A(new_n1312_), .ZN(new_n1499_));
  AND3_X1   g1121(.A1(new_n1494_), .A2(new_n1498_), .A3(new_n1499_), .ZN(new_n1500_));
  AOI21_X1  g1122(.A(new_n1499_), .B1(new_n1494_), .B2(new_n1498_), .ZN(new_n1501_));
  OAI21_X1  g1123(.A(new_n1487_), .B1(new_n1500_), .B2(new_n1501_), .ZN(new_n1502_));
  NAND2_X1  g1124(.A1(new_n1494_), .A2(new_n1498_), .ZN(new_n1503_));
  NAND2_X1  g1125(.A1(new_n1503_), .A2(new_n1312_), .ZN(new_n1504_));
  NAND3_X1  g1126(.A1(new_n1494_), .A2(new_n1498_), .A3(new_n1499_), .ZN(new_n1505_));
  NAND3_X1  g1127(.A1(new_n1504_), .A2(new_n752_), .A3(new_n1505_), .ZN(new_n1506_));
  NAND2_X1  g1128(.A1(new_n1502_), .A2(new_n1506_), .ZN(new_n1507_));
  NAND2_X1  g1129(.A1(new_n1507_), .A2(new_n723_), .ZN(new_n1508_));
  NAND3_X1  g1130(.A1(new_n1502_), .A2(new_n1506_), .A3(new_n722_), .ZN(new_n1509_));
  NAND3_X1  g1131(.A1(new_n1508_), .A2(new_n1328_), .A3(new_n1509_), .ZN(new_n1510_));
  AND3_X1   g1132(.A1(new_n1502_), .A2(new_n1506_), .A3(new_n722_), .ZN(new_n1511_));
  INV_X1    g1133(.A(new_n752_), .ZN(new_n1512_));
  OAI21_X1  g1134(.A(new_n1512_), .B1(new_n1500_), .B2(new_n1501_), .ZN(new_n1513_));
  INV_X1    g1135(.A(KEYINPUT51), .ZN(new_n1514_));
  NAND2_X1  g1136(.A1(new_n1513_), .A2(new_n1514_), .ZN(new_n1515_));
  NAND3_X1  g1137(.A1(new_n1504_), .A2(new_n1066_), .A3(new_n1505_), .ZN(new_n1516_));
  OAI211_X1 g1138(.A(KEYINPUT51), .B(new_n1512_), .C1(new_n1500_), .C2(new_n1501_), .ZN(new_n1517_));
  NAND3_X1  g1139(.A1(new_n1515_), .A2(new_n1516_), .A3(new_n1517_), .ZN(new_n1518_));
  AOI21_X1  g1140(.A(new_n1511_), .B1(new_n1518_), .B2(new_n723_), .ZN(new_n1519_));
  OAI21_X1  g1141(.A(new_n1510_), .B1(new_n1519_), .B2(new_n1328_), .ZN(new_n1520_));
  NAND2_X1  g1142(.A1(new_n1520_), .A2(new_n715_), .ZN(new_n1521_));
  OAI211_X1 g1143(.A(new_n714_), .B(new_n1510_), .C1(new_n1519_), .C2(new_n1328_), .ZN(new_n1522_));
  NAND2_X1  g1144(.A1(new_n1521_), .A2(new_n1522_), .ZN(new_n1523_));
  INV_X1    g1145(.A(new_n1062_), .ZN(new_n1524_));
  NAND2_X1  g1146(.A1(new_n1523_), .A2(new_n1524_), .ZN(new_n1525_));
  AOI211_X1 g1147(.A(new_n791_), .B(new_n1355_), .C1(new_n1062_), .C2(new_n1068_), .ZN(new_n1526_));
  XOR2_X1   g1148(.A(new_n1358_), .B(KEYINPUT52), .Z(new_n1527_));
  AOI211_X1 g1149(.A(new_n537_), .B(new_n1477_), .C1(new_n705_), .C2(new_n780_), .ZN(new_n1528_));
  INV_X1    g1150(.A(new_n539_), .ZN(new_n1529_));
  OAI21_X1  g1151(.A(new_n1068_), .B1(new_n1528_), .B2(new_n1529_), .ZN(new_n1530_));
  AOI21_X1  g1152(.A(new_n1527_), .B1(new_n1530_), .B2(new_n792_), .ZN(new_n1531_));
  NOR2_X1   g1153(.A1(new_n1526_), .A2(new_n1531_), .ZN(new_n1532_));
  AND4_X1   g1154(.A1(new_n745_), .A2(new_n738_), .A3(new_n752_), .A4(new_n756_), .ZN(new_n1533_));
  OAI21_X1  g1155(.A(new_n710_), .B1(new_n1533_), .B2(new_n1311_), .ZN(new_n1534_));
  OAI21_X1  g1156(.A(new_n1309_), .B1(new_n1063_), .B2(new_n1064_), .ZN(new_n1535_));
  NAND3_X1  g1157(.A1(new_n738_), .A2(new_n1307_), .A3(new_n756_), .ZN(new_n1536_));
  NAND2_X1  g1158(.A1(new_n1535_), .A2(new_n1536_), .ZN(new_n1537_));
  INV_X1    g1159(.A(new_n1537_), .ZN(new_n1538_));
  NAND2_X1  g1160(.A1(new_n1534_), .A2(new_n1538_), .ZN(new_n1539_));
  NAND2_X1  g1161(.A1(new_n1320_), .A2(new_n1063_), .ZN(new_n1540_));
  OR2_X1    g1162(.A1(new_n1489_), .A2(new_n1063_), .ZN(new_n1541_));
  INV_X1    g1163(.A(new_n744_), .ZN(new_n1542_));
  AOI21_X1  g1164(.A(new_n1542_), .B1(new_n1488_), .B2(new_n740_), .ZN(new_n1543_));
  NAND3_X1  g1165(.A1(new_n757_), .A2(new_n1543_), .A3(new_n712_), .ZN(new_n1544_));
  NAND3_X1  g1166(.A1(new_n1544_), .A2(new_n1537_), .A3(new_n710_), .ZN(new_n1545_));
  NAND4_X1  g1167(.A1(new_n1539_), .A2(new_n1540_), .A3(new_n1541_), .A4(new_n1545_), .ZN(new_n1546_));
  OAI21_X1  g1168(.A(new_n1540_), .B1(new_n1063_), .B2(new_n1489_), .ZN(new_n1547_));
  AND3_X1   g1169(.A1(new_n1544_), .A2(new_n710_), .A3(new_n1537_), .ZN(new_n1548_));
  AOI21_X1  g1170(.A(new_n1537_), .B1(new_n1544_), .B2(new_n710_), .ZN(new_n1549_));
  OAI21_X1  g1171(.A(new_n1547_), .B1(new_n1548_), .B2(new_n1549_), .ZN(new_n1550_));
  AND3_X1   g1172(.A1(new_n1546_), .A2(new_n1550_), .A3(new_n752_), .ZN(new_n1551_));
  AOI21_X1  g1173(.A(new_n1066_), .B1(new_n1546_), .B2(new_n1550_), .ZN(new_n1552_));
  OAI21_X1  g1174(.A(new_n723_), .B1(new_n1551_), .B2(new_n1552_), .ZN(new_n1553_));
  NOR3_X1   g1175(.A1(new_n1548_), .A2(new_n1549_), .A3(new_n1547_), .ZN(new_n1554_));
  AOI22_X1  g1176(.A1(new_n1539_), .A2(new_n1545_), .B1(new_n1541_), .B2(new_n1540_), .ZN(new_n1555_));
  OAI21_X1  g1177(.A(new_n1487_), .B1(new_n1554_), .B2(new_n1555_), .ZN(new_n1556_));
  NAND3_X1  g1178(.A1(new_n1546_), .A2(new_n1550_), .A3(new_n752_), .ZN(new_n1557_));
  NAND3_X1  g1179(.A1(new_n1556_), .A2(new_n722_), .A3(new_n1557_), .ZN(new_n1558_));
  NAND3_X1  g1180(.A1(new_n1553_), .A2(KEYINPUT49), .A3(new_n1558_), .ZN(new_n1559_));
  INV_X1    g1181(.A(KEYINPUT49), .ZN(new_n1560_));
  OAI211_X1 g1182(.A(new_n1560_), .B(new_n723_), .C1(new_n1551_), .C2(new_n1552_), .ZN(new_n1561_));
  AOI21_X1  g1183(.A(new_n1328_), .B1(new_n1559_), .B2(new_n1561_), .ZN(new_n1562_));
  XNOR2_X1  g1184(.A(new_n1562_), .B(KEYINPUT50), .ZN(new_n1563_));
  OAI21_X1  g1185(.A(new_n752_), .B1(new_n1554_), .B2(new_n1555_), .ZN(new_n1564_));
  NAND3_X1  g1186(.A1(new_n1546_), .A2(new_n1550_), .A3(new_n1487_), .ZN(new_n1565_));
  NAND3_X1  g1187(.A1(new_n1564_), .A2(new_n723_), .A3(new_n1565_), .ZN(new_n1566_));
  NAND2_X1  g1188(.A1(new_n1558_), .A2(new_n1566_), .ZN(new_n1567_));
  NAND2_X1  g1189(.A1(new_n1567_), .A2(new_n1328_), .ZN(new_n1568_));
  AOI21_X1  g1190(.A(new_n714_), .B1(new_n1563_), .B2(new_n1568_), .ZN(new_n1569_));
  AOI21_X1  g1191(.A(new_n1328_), .B1(new_n1558_), .B2(new_n1566_), .ZN(new_n1570_));
  NAND2_X1  g1192(.A1(new_n1559_), .A2(new_n1561_), .ZN(new_n1571_));
  AOI21_X1  g1193(.A(new_n1570_), .B1(new_n1571_), .B2(new_n1328_), .ZN(new_n1572_));
  NOR2_X1   g1194(.A1(new_n1572_), .A2(new_n715_), .ZN(new_n1573_));
  OAI21_X1  g1195(.A(new_n1062_), .B1(new_n1569_), .B2(new_n1573_), .ZN(new_n1574_));
  NAND3_X1  g1196(.A1(new_n1525_), .A2(new_n1532_), .A3(new_n1574_), .ZN(new_n1575_));
  INV_X1    g1197(.A(new_n1355_), .ZN(new_n1576_));
  NAND3_X1  g1198(.A1(new_n1530_), .A2(new_n792_), .A3(new_n1576_), .ZN(new_n1577_));
  OAI21_X1  g1199(.A(new_n1577_), .B1(new_n1069_), .B2(new_n1527_), .ZN(new_n1578_));
  AOI21_X1  g1200(.A(new_n1062_), .B1(new_n1521_), .B2(new_n1522_), .ZN(new_n1579_));
  AOI21_X1  g1201(.A(KEYINPUT53), .B1(new_n1572_), .B2(new_n715_), .ZN(new_n1580_));
  NOR2_X1   g1202(.A1(new_n1580_), .A2(new_n1573_), .ZN(new_n1581_));
  NAND3_X1  g1203(.A1(new_n1572_), .A2(KEYINPUT53), .A3(new_n715_), .ZN(new_n1582_));
  AOI21_X1  g1204(.A(new_n1524_), .B1(new_n1581_), .B2(new_n1582_), .ZN(new_n1583_));
  OAI21_X1  g1205(.A(new_n1578_), .B1(new_n1579_), .B2(new_n1583_), .ZN(new_n1584_));
  AND2_X1   g1206(.A1(new_n1575_), .A2(new_n1584_), .ZN(G338));
  OAI21_X1  g1207(.A(new_n768_), .B1(new_n1375_), .B2(new_n608_), .ZN(new_n1586_));
  XNOR2_X1  g1208(.A(new_n596_), .B(new_n603_), .ZN(new_n1587_));
  XNOR2_X1  g1209(.A(new_n1586_), .B(new_n1587_), .ZN(new_n1588_));
  NOR2_X1   g1210(.A1(new_n772_), .A2(new_n614_), .ZN(new_n1589_));
  XNOR2_X1  g1211(.A(new_n1588_), .B(new_n1589_), .ZN(new_n1590_));
  NAND2_X1  g1212(.A1(new_n776_), .A2(new_n1382_), .ZN(new_n1591_));
  OAI211_X1 g1213(.A(new_n1371_), .B(new_n1591_), .C1(new_n1374_), .C2(new_n621_), .ZN(new_n1592_));
  XNOR2_X1  g1214(.A(new_n1592_), .B(new_n1380_), .ZN(new_n1593_));
  XNOR2_X1  g1215(.A(new_n1590_), .B(new_n1593_), .ZN(new_n1594_));
  NAND2_X1  g1216(.A1(new_n1594_), .A2(new_n1350_), .ZN(new_n1595_));
  INV_X1    g1217(.A(new_n1595_), .ZN(new_n1596_));
  NAND2_X1  g1218(.A1(new_n761_), .A2(new_n575_), .ZN(new_n1597_));
  NAND2_X1  g1219(.A1(new_n567_), .A2(G4427), .ZN(new_n1598_));
  OAI211_X1 g1220(.A(new_n1406_), .B(new_n1597_), .C1(new_n575_), .C2(new_n1598_), .ZN(new_n1599_));
  INV_X1    g1221(.A(new_n576_), .ZN(new_n1600_));
  NAND4_X1  g1222(.A1(new_n1600_), .A2(G4427), .A3(new_n567_), .A4(new_n574_), .ZN(new_n1601_));
  AND2_X1   g1223(.A1(new_n1599_), .A2(new_n1601_), .ZN(new_n1602_));
  NAND3_X1  g1224(.A1(new_n1602_), .A2(new_n1396_), .A3(new_n760_), .ZN(new_n1603_));
  INV_X1    g1225(.A(new_n1603_), .ZN(new_n1604_));
  AOI21_X1  g1226(.A(new_n1602_), .B1(new_n1396_), .B2(new_n760_), .ZN(new_n1605_));
  NOR3_X1   g1227(.A1(new_n1604_), .A2(new_n1605_), .A3(new_n571_), .ZN(new_n1606_));
  NAND2_X1  g1228(.A1(new_n1599_), .A2(new_n1601_), .ZN(new_n1607_));
  NAND2_X1  g1229(.A1(new_n1397_), .A2(new_n1607_), .ZN(new_n1608_));
  AOI22_X1  g1230(.A1(new_n1608_), .A2(new_n1603_), .B1(new_n570_), .B2(new_n564_), .ZN(new_n1609_));
  NOR2_X1   g1231(.A1(new_n1606_), .A2(new_n1609_), .ZN(new_n1610_));
  INV_X1    g1232(.A(new_n1610_), .ZN(new_n1611_));
  OAI21_X1  g1233(.A(new_n571_), .B1(new_n1604_), .B2(new_n1605_), .ZN(new_n1612_));
  INV_X1    g1234(.A(KEYINPUT58), .ZN(new_n1613_));
  NAND2_X1  g1235(.A1(new_n1612_), .A2(new_n1613_), .ZN(new_n1614_));
  AOI21_X1  g1236(.A(new_n1402_), .B1(new_n1614_), .B2(new_n1390_), .ZN(new_n1615_));
  AOI211_X1 g1237(.A(new_n581_), .B(new_n588_), .C1(new_n1612_), .C2(new_n1613_), .ZN(new_n1616_));
  OAI21_X1  g1238(.A(new_n1611_), .B1(new_n1615_), .B2(new_n1616_), .ZN(new_n1617_));
  OAI21_X1  g1239(.A(new_n1390_), .B1(new_n1609_), .B2(KEYINPUT58), .ZN(new_n1618_));
  NAND2_X1  g1240(.A1(new_n1618_), .A2(new_n588_), .ZN(new_n1619_));
  NAND3_X1  g1241(.A1(new_n1614_), .A2(new_n1390_), .A3(new_n1402_), .ZN(new_n1620_));
  NAND3_X1  g1242(.A1(new_n1619_), .A2(new_n1620_), .A3(new_n1610_), .ZN(new_n1621_));
  NAND3_X1  g1243(.A1(new_n1617_), .A2(new_n1621_), .A3(new_n779_), .ZN(new_n1622_));
  NAND2_X1  g1244(.A1(new_n1622_), .A2(new_n1350_), .ZN(new_n1623_));
  NAND2_X1  g1245(.A1(new_n778_), .A2(new_n625_), .ZN(new_n1624_));
  NAND2_X1  g1246(.A1(new_n1623_), .A2(new_n1624_), .ZN(new_n1625_));
  OAI21_X1  g1247(.A(new_n585_), .B1(new_n762_), .B2(new_n587_), .ZN(new_n1626_));
  NAND2_X1  g1248(.A1(new_n1598_), .A2(new_n576_), .ZN(new_n1627_));
  XNOR2_X1  g1249(.A(new_n761_), .B(new_n575_), .ZN(new_n1628_));
  OAI21_X1  g1250(.A(new_n1627_), .B1(new_n1628_), .B2(new_n576_), .ZN(new_n1629_));
  XNOR2_X1  g1251(.A(new_n1626_), .B(new_n1629_), .ZN(new_n1630_));
  XNOR2_X1  g1252(.A(new_n571_), .B(new_n1390_), .ZN(new_n1631_));
  XNOR2_X1  g1253(.A(new_n1630_), .B(new_n1631_), .ZN(new_n1632_));
  NAND2_X1  g1254(.A1(new_n1625_), .A2(new_n1632_), .ZN(new_n1633_));
  NAND2_X1  g1255(.A1(new_n1617_), .A2(new_n1621_), .ZN(new_n1634_));
  NAND2_X1  g1256(.A1(new_n1634_), .A2(new_n1389_), .ZN(new_n1635_));
  AOI21_X1  g1257(.A(new_n1596_), .B1(new_n1633_), .B2(new_n1635_), .ZN(new_n1636_));
  INV_X1    g1258(.A(KEYINPUT54), .ZN(new_n1637_));
  AOI21_X1  g1259(.A(new_n615_), .B1(new_n622_), .B2(new_n1637_), .ZN(new_n1638_));
  NAND2_X1  g1260(.A1(new_n1373_), .A2(new_n1638_), .ZN(new_n1639_));
  NAND3_X1  g1261(.A1(new_n622_), .A2(new_n1637_), .A3(new_n613_), .ZN(new_n1640_));
  NAND2_X1  g1262(.A1(new_n1639_), .A2(new_n1640_), .ZN(new_n1641_));
  NAND2_X1  g1263(.A1(new_n1374_), .A2(new_n607_), .ZN(new_n1642_));
  AOI21_X1  g1264(.A(new_n1641_), .B1(new_n1642_), .B2(new_n768_), .ZN(new_n1643_));
  INV_X1    g1265(.A(new_n1643_), .ZN(new_n1644_));
  NAND3_X1  g1266(.A1(new_n1642_), .A2(new_n768_), .A3(new_n1641_), .ZN(new_n1645_));
  NAND3_X1  g1267(.A1(new_n1644_), .A2(new_n623_), .A3(new_n1645_), .ZN(new_n1646_));
  AND3_X1   g1268(.A1(new_n1642_), .A2(new_n768_), .A3(new_n1641_), .ZN(new_n1647_));
  OAI21_X1  g1269(.A(new_n624_), .B1(new_n1647_), .B2(new_n1643_), .ZN(new_n1648_));
  NAND2_X1  g1270(.A1(new_n1646_), .A2(new_n1648_), .ZN(new_n1649_));
  NAND2_X1  g1271(.A1(new_n1649_), .A2(new_n1374_), .ZN(new_n1650_));
  INV_X1    g1272(.A(new_n1374_), .ZN(new_n1651_));
  NAND3_X1  g1273(.A1(new_n1646_), .A2(new_n1648_), .A3(new_n1651_), .ZN(new_n1652_));
  AOI21_X1  g1274(.A(new_n616_), .B1(new_n1650_), .B2(new_n1652_), .ZN(new_n1653_));
  NOR3_X1   g1275(.A1(new_n1653_), .A2(KEYINPUT55), .A3(new_n1378_), .ZN(new_n1654_));
  AND3_X1   g1276(.A1(new_n1646_), .A2(new_n1651_), .A3(new_n1648_), .ZN(new_n1655_));
  AOI21_X1  g1277(.A(new_n1651_), .B1(new_n1646_), .B2(new_n1648_), .ZN(new_n1656_));
  NOR3_X1   g1278(.A1(new_n1655_), .A2(new_n1656_), .A3(new_n771_), .ZN(new_n1657_));
  OAI21_X1  g1279(.A(new_n1378_), .B1(new_n1657_), .B2(new_n1653_), .ZN(new_n1658_));
  OAI21_X1  g1280(.A(new_n771_), .B1(new_n1655_), .B2(new_n1656_), .ZN(new_n1659_));
  NAND3_X1  g1281(.A1(new_n1650_), .A2(new_n616_), .A3(new_n1652_), .ZN(new_n1660_));
  NAND3_X1  g1282(.A1(new_n1659_), .A2(new_n1660_), .A3(new_n596_), .ZN(new_n1661_));
  AOI21_X1  g1283(.A(new_n1654_), .B1(new_n1658_), .B2(new_n1661_), .ZN(new_n1662_));
  NOR4_X1   g1284(.A1(new_n1653_), .A2(new_n1660_), .A3(KEYINPUT55), .A4(new_n1378_), .ZN(new_n1663_));
  OAI21_X1  g1285(.A(new_n1385_), .B1(new_n1662_), .B2(new_n1663_), .ZN(new_n1664_));
  NAND3_X1  g1286(.A1(new_n1658_), .A2(new_n603_), .A3(new_n1661_), .ZN(new_n1665_));
  NAND2_X1  g1287(.A1(new_n1665_), .A2(KEYINPUT56), .ZN(new_n1666_));
  INV_X1    g1288(.A(KEYINPUT56), .ZN(new_n1667_));
  NAND4_X1  g1289(.A1(new_n1658_), .A2(new_n1667_), .A3(new_n603_), .A4(new_n1661_), .ZN(new_n1668_));
  NAND4_X1  g1290(.A1(new_n1664_), .A2(new_n610_), .A3(new_n1666_), .A4(new_n1668_), .ZN(new_n1669_));
  INV_X1    g1291(.A(KEYINPUT57), .ZN(new_n1670_));
  NAND2_X1  g1292(.A1(new_n1669_), .A2(new_n1670_), .ZN(new_n1671_));
  NAND2_X1  g1293(.A1(new_n1666_), .A2(new_n1668_), .ZN(new_n1672_));
  INV_X1    g1294(.A(new_n1672_), .ZN(new_n1673_));
  NAND4_X1  g1295(.A1(new_n1673_), .A2(KEYINPUT57), .A3(new_n610_), .A4(new_n1664_), .ZN(new_n1674_));
  OAI21_X1  g1296(.A(new_n603_), .B1(new_n1662_), .B2(new_n1663_), .ZN(new_n1675_));
  NAND3_X1  g1297(.A1(new_n1658_), .A2(new_n1385_), .A3(new_n1661_), .ZN(new_n1676_));
  NAND3_X1  g1298(.A1(new_n1675_), .A2(new_n1380_), .A3(new_n1676_), .ZN(new_n1677_));
  NAND3_X1  g1299(.A1(new_n1671_), .A2(new_n1674_), .A3(new_n1677_), .ZN(new_n1678_));
  NAND2_X1  g1300(.A1(new_n1678_), .A2(new_n1369_), .ZN(new_n1679_));
  INV_X1    g1301(.A(KEYINPUT55), .ZN(new_n1680_));
  NAND3_X1  g1302(.A1(new_n1659_), .A2(new_n1680_), .A3(new_n596_), .ZN(new_n1681_));
  AND3_X1   g1303(.A1(new_n1659_), .A2(new_n1660_), .A3(new_n596_), .ZN(new_n1682_));
  AOI21_X1  g1304(.A(new_n596_), .B1(new_n1659_), .B2(new_n1660_), .ZN(new_n1683_));
  OAI21_X1  g1305(.A(new_n1681_), .B1(new_n1682_), .B2(new_n1683_), .ZN(new_n1684_));
  NAND3_X1  g1306(.A1(new_n1658_), .A2(new_n1654_), .A3(new_n1661_), .ZN(new_n1685_));
  AOI21_X1  g1307(.A(new_n603_), .B1(new_n1684_), .B2(new_n1685_), .ZN(new_n1686_));
  OAI21_X1  g1308(.A(new_n1380_), .B1(new_n1672_), .B2(new_n1686_), .ZN(new_n1687_));
  AND2_X1   g1309(.A1(new_n1687_), .A2(new_n1669_), .ZN(new_n1688_));
  OAI21_X1  g1310(.A(new_n1595_), .B1(new_n1688_), .B2(new_n1350_), .ZN(new_n1689_));
  AOI22_X1  g1311(.A1(new_n1625_), .A2(new_n1632_), .B1(new_n1634_), .B2(new_n1389_), .ZN(new_n1690_));
  AOI22_X1  g1312(.A1(new_n1636_), .A2(new_n1679_), .B1(new_n1689_), .B2(new_n1690_), .ZN(G370));
  OAI21_X1  g1313(.A(new_n671_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n1692_));
  NAND2_X1  g1314(.A1(new_n657_), .A2(new_n439_), .ZN(new_n1693_));
  NAND2_X1  g1315(.A1(new_n1692_), .A2(new_n1693_), .ZN(new_n1694_));
  OAI211_X1 g1316(.A(new_n1075_), .B(new_n1694_), .C1(new_n438_), .C2(new_n1078_), .ZN(new_n1695_));
  OAI211_X1 g1317(.A(new_n651_), .B(new_n1074_), .C1(new_n1078_), .C2(new_n438_), .ZN(new_n1696_));
  NAND3_X1  g1318(.A1(new_n1696_), .A2(new_n1693_), .A3(new_n1692_), .ZN(new_n1697_));
  NAND2_X1  g1319(.A1(new_n1695_), .A2(new_n1697_), .ZN(new_n1698_));
  NAND2_X1  g1320(.A1(new_n1085_), .A2(new_n1079_), .ZN(new_n1699_));
  INV_X1    g1321(.A(KEYINPUT59), .ZN(new_n1700_));
  NAND2_X1  g1322(.A1(new_n1699_), .A2(new_n1700_), .ZN(new_n1701_));
  NAND2_X1  g1323(.A1(new_n1084_), .A2(new_n438_), .ZN(new_n1702_));
  NAND3_X1  g1324(.A1(new_n1085_), .A2(KEYINPUT59), .A3(new_n1079_), .ZN(new_n1703_));
  NAND3_X1  g1325(.A1(new_n1701_), .A2(new_n1702_), .A3(new_n1703_), .ZN(new_n1704_));
  NAND2_X1  g1326(.A1(new_n1698_), .A2(new_n1704_), .ZN(new_n1705_));
  AND2_X1   g1327(.A1(new_n1701_), .A2(new_n1703_), .ZN(new_n1706_));
  NAND4_X1  g1328(.A1(new_n1706_), .A2(new_n1697_), .A3(new_n1702_), .A4(new_n1695_), .ZN(new_n1707_));
  NAND2_X1  g1329(.A1(new_n1705_), .A2(new_n1707_), .ZN(new_n1708_));
  NAND2_X1  g1330(.A1(new_n1708_), .A2(new_n662_), .ZN(new_n1709_));
  NAND3_X1  g1331(.A1(new_n1705_), .A2(new_n1707_), .A3(new_n1077_), .ZN(new_n1710_));
  NAND3_X1  g1332(.A1(new_n1709_), .A2(KEYINPUT60), .A3(new_n1710_), .ZN(new_n1711_));
  OR2_X1    g1333(.A1(new_n1710_), .A2(KEYINPUT60), .ZN(new_n1712_));
  AOI21_X1  g1334(.A(new_n1082_), .B1(new_n1711_), .B2(new_n1712_), .ZN(new_n1713_));
  AOI21_X1  g1335(.A(new_n664_), .B1(new_n1709_), .B2(new_n1710_), .ZN(new_n1714_));
  OAI21_X1  g1336(.A(new_n646_), .B1(new_n1713_), .B2(new_n1714_), .ZN(new_n1715_));
  INV_X1    g1337(.A(KEYINPUT61), .ZN(new_n1716_));
  NAND2_X1  g1338(.A1(new_n1715_), .A2(new_n1716_), .ZN(new_n1717_));
  NAND2_X1  g1339(.A1(new_n1711_), .A2(new_n1712_), .ZN(new_n1718_));
  NAND2_X1  g1340(.A1(new_n1718_), .A2(new_n664_), .ZN(new_n1719_));
  NAND3_X1  g1341(.A1(new_n1711_), .A2(new_n1712_), .A3(new_n1082_), .ZN(new_n1720_));
  NAND3_X1  g1342(.A1(new_n1719_), .A2(new_n1090_), .A3(new_n1720_), .ZN(new_n1721_));
  OAI211_X1 g1343(.A(KEYINPUT61), .B(new_n646_), .C1(new_n1713_), .C2(new_n1714_), .ZN(new_n1722_));
  NAND3_X1  g1344(.A1(new_n1717_), .A2(new_n1721_), .A3(new_n1722_), .ZN(new_n1723_));
  NAND2_X1  g1345(.A1(new_n1723_), .A2(new_n653_), .ZN(new_n1724_));
  INV_X1    g1346(.A(new_n1720_), .ZN(new_n1725_));
  OAI21_X1  g1347(.A(new_n1091_), .B1(new_n1725_), .B2(new_n1713_), .ZN(new_n1726_));
  INV_X1    g1348(.A(new_n1714_), .ZN(new_n1727_));
  NAND3_X1  g1349(.A1(new_n1719_), .A2(new_n1073_), .A3(new_n1727_), .ZN(new_n1728_));
  AND3_X1   g1350(.A1(new_n1726_), .A2(new_n1728_), .A3(new_n1076_), .ZN(new_n1729_));
  INV_X1    g1351(.A(new_n1729_), .ZN(new_n1730_));
  NAND2_X1  g1352(.A1(new_n1724_), .A2(new_n1730_), .ZN(new_n1731_));
  NAND2_X1  g1353(.A1(new_n1731_), .A2(G4526), .ZN(new_n1732_));
  AOI21_X1  g1354(.A(new_n1096_), .B1(new_n692_), .B2(new_n686_), .ZN(new_n1733_));
  INV_X1    g1355(.A(KEYINPUT63), .ZN(new_n1734_));
  AOI21_X1  g1356(.A(new_n1097_), .B1(new_n1733_), .B2(new_n1734_), .ZN(new_n1735_));
  XNOR2_X1  g1357(.A(new_n1735_), .B(new_n680_), .ZN(new_n1736_));
  NOR2_X1   g1358(.A1(new_n1733_), .A2(new_n1734_), .ZN(new_n1737_));
  XNOR2_X1  g1359(.A(new_n1737_), .B(new_n1100_), .ZN(new_n1738_));
  OR2_X1    g1360(.A1(new_n1736_), .A2(new_n1738_), .ZN(new_n1739_));
  NAND2_X1  g1361(.A1(new_n1736_), .A2(new_n1738_), .ZN(new_n1740_));
  NAND2_X1  g1362(.A1(new_n1739_), .A2(new_n1740_), .ZN(new_n1741_));
  NOR2_X1   g1363(.A1(new_n1741_), .A2(new_n688_), .ZN(new_n1742_));
  NAND2_X1  g1364(.A1(new_n1741_), .A2(new_n688_), .ZN(new_n1743_));
  INV_X1    g1365(.A(new_n1743_), .ZN(new_n1744_));
  OAI22_X1  g1366(.A1(new_n1742_), .A2(new_n1744_), .B1(new_n694_), .B2(new_n693_), .ZN(new_n1745_));
  INV_X1    g1367(.A(new_n1742_), .ZN(new_n1746_));
  NAND3_X1  g1368(.A1(new_n1746_), .A2(new_n695_), .A3(new_n1743_), .ZN(new_n1747_));
  NAND2_X1  g1369(.A1(new_n1745_), .A2(new_n1747_), .ZN(new_n1748_));
  OAI21_X1  g1370(.A(new_n638_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n1749_));
  NAND2_X1  g1371(.A1(new_n1748_), .A2(new_n1749_), .ZN(new_n1750_));
  OAI21_X1  g1372(.A(new_n699_), .B1(new_n698_), .B2(new_n693_), .ZN(new_n1751_));
  XNOR2_X1  g1373(.A(new_n1751_), .B(new_n680_), .ZN(new_n1752_));
  XNOR2_X1  g1374(.A(new_n1752_), .B(new_n688_), .ZN(new_n1753_));
  INV_X1    g1375(.A(new_n1753_), .ZN(new_n1754_));
  XNOR2_X1  g1376(.A(new_n1100_), .B(new_n695_), .ZN(new_n1755_));
  XOR2_X1   g1377(.A(new_n702_), .B(new_n1755_), .Z(new_n1756_));
  OR2_X1    g1378(.A1(new_n1754_), .A2(new_n1756_), .ZN(new_n1757_));
  AOI22_X1  g1379(.A1(new_n1754_), .A2(new_n1756_), .B1(G4526), .B2(new_n675_), .ZN(new_n1758_));
  NAND3_X1  g1380(.A1(new_n1750_), .A2(new_n1757_), .A3(new_n1758_), .ZN(new_n1759_));
  NAND3_X1  g1381(.A1(new_n1745_), .A2(new_n675_), .A3(new_n1747_), .ZN(new_n1760_));
  NAND2_X1  g1382(.A1(new_n1759_), .A2(new_n1760_), .ZN(new_n1761_));
  NAND2_X1  g1383(.A1(new_n672_), .A2(new_n652_), .ZN(new_n1762_));
  NAND2_X1  g1384(.A1(new_n1762_), .A2(new_n1077_), .ZN(new_n1763_));
  NAND3_X1  g1385(.A1(new_n672_), .A2(new_n652_), .A3(new_n662_), .ZN(new_n1764_));
  INV_X1    g1386(.A(new_n436_), .ZN(new_n1765_));
  NAND2_X1  g1387(.A1(new_n1092_), .A2(new_n667_), .ZN(new_n1766_));
  AOI21_X1  g1388(.A(new_n1765_), .B1(new_n1766_), .B2(new_n644_), .ZN(new_n1767_));
  NOR2_X1   g1389(.A1(new_n1084_), .A2(new_n436_), .ZN(new_n1768_));
  NOR2_X1   g1390(.A1(new_n1767_), .A2(new_n1768_), .ZN(new_n1769_));
  INV_X1    g1391(.A(new_n1769_), .ZN(new_n1770_));
  AND3_X1   g1392(.A1(new_n1763_), .A2(new_n1764_), .A3(new_n1770_), .ZN(new_n1771_));
  AOI21_X1  g1393(.A(new_n1770_), .B1(new_n1763_), .B2(new_n1764_), .ZN(new_n1772_));
  XNOR2_X1  g1394(.A(new_n671_), .B(new_n439_), .ZN(new_n1773_));
  INV_X1    g1395(.A(new_n1773_), .ZN(new_n1774_));
  OR3_X1    g1396(.A1(new_n1771_), .A2(new_n1772_), .A3(new_n1774_), .ZN(new_n1775_));
  INV_X1    g1397(.A(KEYINPUT62), .ZN(new_n1776_));
  OAI21_X1  g1398(.A(new_n1774_), .B1(new_n1771_), .B2(new_n1772_), .ZN(new_n1777_));
  NAND4_X1  g1399(.A1(new_n1775_), .A2(new_n1776_), .A3(new_n1082_), .A4(new_n1777_), .ZN(new_n1778_));
  NAND2_X1  g1400(.A1(new_n1778_), .A2(new_n1091_), .ZN(new_n1779_));
  AOI21_X1  g1401(.A(new_n1082_), .B1(new_n1775_), .B2(new_n1777_), .ZN(new_n1780_));
  NOR2_X1   g1402(.A1(new_n1780_), .A2(new_n1776_), .ZN(new_n1781_));
  NAND3_X1  g1403(.A1(new_n1775_), .A2(new_n1082_), .A3(new_n1777_), .ZN(new_n1782_));
  AOI21_X1  g1404(.A(new_n1779_), .B1(new_n1781_), .B2(new_n1782_), .ZN(new_n1783_));
  INV_X1    g1405(.A(new_n1782_), .ZN(new_n1784_));
  NOR3_X1   g1406(.A1(new_n1784_), .A2(new_n646_), .A3(new_n1780_), .ZN(new_n1785_));
  OR3_X1    g1407(.A1(new_n1783_), .A2(new_n1785_), .A3(new_n653_), .ZN(new_n1786_));
  OAI21_X1  g1408(.A(new_n653_), .B1(new_n1783_), .B2(new_n1785_), .ZN(new_n1787_));
  NAND3_X1  g1409(.A1(new_n1786_), .A2(new_n1787_), .A3(new_n440_), .ZN(new_n1788_));
  AND2_X1   g1410(.A1(new_n1761_), .A2(new_n1788_), .ZN(new_n1789_));
  AOI21_X1  g1411(.A(new_n1076_), .B1(new_n1726_), .B2(new_n1728_), .ZN(new_n1790_));
  OAI21_X1  g1412(.A(G4526), .B1(new_n1729_), .B2(new_n1790_), .ZN(new_n1791_));
  NAND2_X1  g1413(.A1(new_n1791_), .A2(new_n1788_), .ZN(new_n1792_));
  INV_X1    g1414(.A(new_n1761_), .ZN(new_n1793_));
  AOI22_X1  g1415(.A1(new_n1732_), .A2(new_n1789_), .B1(new_n1792_), .B2(new_n1793_), .ZN(G399));
endmodule


