//Secret key is'0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_c7552" written by ABC on Sun Nov 20 19:50:25 2022

module locked_c7552 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G5, G9, G12, G15, G18, G23, G26, G29,
    G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59,
    G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77,
    G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97,
    G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121,
    G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151,
    G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163,
    G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175,
    G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187,
    G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199,
    G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211,
    G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223,
    G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235,
    G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469,
    G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230,
    G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717,
    G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410,
    G4415, G4420, G4427, G4432, G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G5, G9, G12, G15, G18, G23,
    G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57,
    G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75,
    G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89,
    G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115,
    G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147,
    G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161,
    G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173,
    G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185,
    G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197,
    G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209,
    G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221,
    G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233,
    G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459,
    G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218,
    G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705,
    G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400,
    G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_n484_, new_n491_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1263_, new_n1265_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1462_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1505_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1535_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1561_, new_n1563_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1612_, new_n1613_, new_n1614_, new_n1616_, new_n1617_,
    new_n1618_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_;
  BUF_X1    g0000(.A(G1), .Z(G2));
  BUF_X1    g0001(.A(G1), .Z(G3));
  XOR2_X1   g0002(.A(KEYINPUT0), .B(G1459), .Z(G450));
  BUF_X1    g0003(.A(G1469), .Z(G448));
  BUF_X1    g0004(.A(G1480), .Z(G444));
  BUF_X1    g0005(.A(G1486), .Z(G442));
  BUF_X1    g0006(.A(G1492), .Z(G440));
  BUF_X1    g0007(.A(G1496), .Z(G438));
  BUF_X1    g0008(.A(G2208), .Z(G496));
  BUF_X1    g0009(.A(G2218), .Z(G494));
  BUF_X1    g0010(.A(G2224), .Z(G492));
  BUF_X1    g0011(.A(G2230), .Z(G490));
  BUF_X1    g0012(.A(G2236), .Z(G488));
  BUF_X1    g0013(.A(G2239), .Z(G486));
  BUF_X1    g0014(.A(G2247), .Z(G484));
  BUF_X1    g0015(.A(G2253), .Z(G482));
  BUF_X1    g0016(.A(G2256), .Z(G480));
  BUF_X1    g0017(.A(G3698), .Z(G560));
  BUF_X1    g0018(.A(G3701), .Z(G542));
  BUF_X1    g0019(.A(G3705), .Z(G558));
  BUF_X1    g0020(.A(G3711), .Z(G556));
  BUF_X1    g0021(.A(G3717), .Z(G554));
  BUF_X1    g0022(.A(G3723), .Z(G552));
  BUF_X1    g0023(.A(G3729), .Z(G550));
  BUF_X1    g0024(.A(G3737), .Z(G548));
  BUF_X1    g0025(.A(G3743), .Z(G546));
  BUF_X1    g0026(.A(G3749), .Z(G544));
  BUF_X1    g0027(.A(G4393), .Z(G540));
  BUF_X1    g0028(.A(G4400), .Z(G538));
  BUF_X1    g0029(.A(G4405), .Z(G536));
  BUF_X1    g0030(.A(G4410), .Z(G534));
  BUF_X1    g0031(.A(G4415), .Z(G532));
  BUF_X1    g0032(.A(G4420), .Z(G530));
  BUF_X1    g0033(.A(G4427), .Z(G528));
  XNOR2_X1  g0034(.A(KEYINPUT1), .B(G4432), .ZN(G526));
  BUF_X1    g0035(.A(G4437), .Z(G524));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G15), .ZN(G279));
  BUF_X1    g0037(.A(G1462), .Z(G436));
  BUF_X1    g0038(.A(G2211), .Z(G478));
  BUF_X1    g0039(.A(G4394), .Z(G522));
  OR2_X1    g0040(.A1(G5), .A2(G57), .ZN(G402));
  NAND4_X1  g0041(.A1(G150), .A2(G184), .A3(G228), .A4(G240), .ZN(new_n484_));
  XOR2_X1   g0042(.A(new_n484_), .B(KEYINPUT3), .Z(G404));
  NAND4_X1  g0043(.A1(G152), .A2(G210), .A3(G218), .A4(G230), .ZN(G406));
  NAND4_X1  g0044(.A1(G182), .A2(G183), .A3(G185), .A4(G186), .ZN(G408));
  NAND4_X1  g0045(.A1(G162), .A2(G172), .A3(G188), .A4(G199), .ZN(G410));
  BUF_X1    g0046(.A(G1), .Z(G432));
  BUF_X1    g0047(.A(G106), .Z(G446));
  INV_X1    g0048(.A(G5), .ZN(new_n491_));
  NAND2_X1  g0049(.A1(new_n491_), .A2(G1197), .ZN(G284));
  INV_X1    g0050(.A(G15), .ZN(G286));
  NAND2_X1  g0051(.A1(new_n491_), .A2(G1197), .ZN(G289));
  NAND3_X1  g0052(.A1(new_n491_), .A2(G133), .A3(G134), .ZN(G292));
  INV_X1    g0053(.A(G15), .ZN(G341));
  NAND3_X1  g0054(.A1(new_n491_), .A2(G133), .A3(G134), .ZN(G281));
  BUF_X1    g0055(.A(G1), .Z(G453));
  AND2_X1   g0056(.A1(G1), .A2(G163), .ZN(G278));
  INV_X1    g0057(.A(G41), .ZN(new_n500_));
  NOR3_X1   g0058(.A1(new_n500_), .A2(G18), .A3(G3701), .ZN(new_n501_));
  INV_X1    g0059(.A(G3701), .ZN(new_n502_));
  NOR3_X1   g0060(.A1(new_n502_), .A2(G18), .A3(G41), .ZN(new_n503_));
  NOR2_X1   g0061(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g0062(.A(G4526), .ZN(new_n505_));
  XNOR2_X1  g0063(.A(new_n504_), .B(new_n505_), .ZN(G373));
  INV_X1    g0064(.A(G18), .ZN(new_n507_));
  OR2_X1    g0065(.A1(new_n507_), .A2(G157), .ZN(new_n508_));
  NAND2_X1  g0066(.A1(G9), .A2(G12), .ZN(new_n509_));
  NAND2_X1  g0067(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g0068(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g0069(.A(G2236), .ZN(new_n512_));
  NAND2_X1  g0070(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g0071(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g0072(.A1(G18), .A2(G160), .ZN(new_n515_));
  INV_X1    g0073(.A(G138), .ZN(new_n516_));
  OAI21_X1  g0074(.A(new_n515_), .B1(new_n516_), .B2(G18), .ZN(new_n517_));
  INV_X1    g0075(.A(G2218), .ZN(new_n518_));
  NAND2_X1  g0076(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g0077(.A(KEYINPUT20), .ZN(new_n520_));
  NAND2_X1  g0078(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g0079(.A1(new_n507_), .A2(G144), .ZN(new_n522_));
  NAND2_X1  g0080(.A1(G18), .A2(G159), .ZN(new_n523_));
  NAND2_X1  g0081(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g0082(.A(G2224), .ZN(new_n525_));
  NAND2_X1  g0083(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g0084(.A1(new_n517_), .A2(KEYINPUT20), .A3(new_n518_), .ZN(new_n527_));
  NAND3_X1  g0085(.A1(new_n521_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g0086(.A(G144), .ZN(new_n529_));
  OAI211_X1 g0087(.A(new_n523_), .B(G2224), .C1(G18), .C2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g0088(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g0089(.A(new_n515_), .B(G2218), .C1(G18), .C2(new_n516_), .ZN(new_n532_));
  AND2_X1   g0090(.A1(new_n519_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g0091(.A(G147), .ZN(new_n534_));
  OAI21_X1  g0092(.A(KEYINPUT10), .B1(new_n534_), .B2(G18), .ZN(new_n535_));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n536_));
  NAND3_X1  g0094(.A1(new_n536_), .A2(new_n507_), .A3(G147), .ZN(new_n537_));
  NAND2_X1  g0095(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g0096(.A1(G18), .A2(G151), .ZN(new_n539_));
  AOI21_X1  g0097(.A(G2211), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g0098(.A(new_n530_), .ZN(new_n541_));
  AOI21_X1  g0099(.A(G2224), .B1(new_n522_), .B2(new_n523_), .ZN(new_n542_));
  NOR2_X1   g0100(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g0101(.A1(new_n533_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g0102(.A1(new_n531_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g0103(.A(G2230), .ZN(new_n546_));
  NAND2_X1  g0104(.A1(G18), .A2(G158), .ZN(new_n547_));
  INV_X1    g0105(.A(G135), .ZN(new_n548_));
  OAI21_X1  g0106(.A(new_n547_), .B1(new_n548_), .B2(G18), .ZN(new_n549_));
  INV_X1    g0107(.A(KEYINPUT8), .ZN(new_n550_));
  NAND2_X1  g0108(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g0109(.A(new_n547_), .B(KEYINPUT8), .C1(G18), .C2(new_n548_), .ZN(new_n552_));
  AOI21_X1  g0110(.A(new_n546_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g0111(.A(new_n547_), .B(new_n546_), .C1(G18), .C2(new_n548_), .ZN(new_n554_));
  NAND2_X1  g0112(.A1(new_n554_), .A2(KEYINPUT9), .ZN(new_n555_));
  NAND2_X1  g0113(.A1(new_n507_), .A2(G135), .ZN(new_n556_));
  INV_X1    g0114(.A(KEYINPUT9), .ZN(new_n557_));
  NAND4_X1  g0115(.A1(new_n556_), .A2(new_n557_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n558_));
  NAND2_X1  g0116(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g0117(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g0118(.A1(new_n511_), .A2(new_n512_), .ZN(new_n561_));
  NOR2_X1   g0119(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g0120(.A(new_n514_), .B1(new_n545_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g0121(.A(KEYINPUT21), .ZN(new_n564_));
  OR2_X1    g0122(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g0123(.A1(new_n514_), .A2(new_n561_), .ZN(new_n566_));
  NAND2_X1  g0124(.A1(new_n551_), .A2(new_n552_), .ZN(new_n567_));
  NAND2_X1  g0125(.A1(new_n567_), .A2(new_n546_), .ZN(new_n568_));
  INV_X1    g0126(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g0127(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g0128(.A1(new_n563_), .A2(new_n564_), .ZN(new_n571_));
  NAND3_X1  g0129(.A1(new_n565_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AND2_X1   g0130(.A1(G9), .A2(G12), .ZN(new_n573_));
  INV_X1    g0131(.A(G154), .ZN(new_n574_));
  AOI21_X1  g0132(.A(new_n573_), .B1(G18), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g0133(.A(G2253), .ZN(new_n576_));
  NOR2_X1   g0134(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g0135(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g0136(.A1(new_n575_), .A2(new_n576_), .ZN(new_n579_));
  NAND2_X1  g0137(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g0138(.A(new_n580_), .B(KEYINPUT5), .ZN(new_n581_));
  OAI21_X1  g0139(.A(new_n509_), .B1(new_n507_), .B2(G155), .ZN(new_n582_));
  OR2_X1    g0140(.A1(new_n582_), .A2(KEYINPUT6), .ZN(new_n583_));
  NAND2_X1  g0141(.A1(new_n582_), .A2(KEYINPUT6), .ZN(new_n584_));
  NAND3_X1  g0142(.A1(new_n583_), .A2(G2247), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g0143(.A(new_n582_), .ZN(new_n586_));
  INV_X1    g0144(.A(G2247), .ZN(new_n587_));
  NAND2_X1  g0145(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g0146(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g0147(.A(G156), .ZN(new_n590_));
  NAND2_X1  g0148(.A1(new_n590_), .A2(G18), .ZN(new_n591_));
  NAND2_X1  g0149(.A1(new_n591_), .A2(new_n509_), .ZN(new_n592_));
  NAND2_X1  g0150(.A1(new_n592_), .A2(G2239), .ZN(new_n593_));
  INV_X1    g0151(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g0152(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g0153(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g0154(.A(new_n592_), .ZN(new_n597_));
  INV_X1    g0155(.A(G2239), .ZN(new_n598_));
  NAND2_X1  g0156(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g0157(.A(new_n599_), .ZN(new_n600_));
  OAI21_X1  g0158(.A(new_n509_), .B1(new_n507_), .B2(G153), .ZN(new_n601_));
  XNOR2_X1  g0159(.A(new_n601_), .B(KEYINPUT7), .ZN(new_n602_));
  OR2_X1    g0160(.A1(new_n602_), .A2(G2256), .ZN(new_n603_));
  NAND2_X1  g0161(.A1(new_n602_), .A2(G2256), .ZN(new_n604_));
  NAND2_X1  g0162(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR4_X1   g0163(.A1(new_n581_), .A2(new_n596_), .A3(new_n600_), .A4(new_n605_), .ZN(new_n606_));
  NAND2_X1  g0164(.A1(new_n572_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g0165(.A1(new_n583_), .A2(new_n584_), .ZN(new_n608_));
  NAND2_X1  g0166(.A1(new_n608_), .A2(new_n587_), .ZN(new_n609_));
  NAND2_X1  g0167(.A1(new_n609_), .A2(new_n579_), .ZN(new_n610_));
  INV_X1    g0168(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g0169(.A1(new_n585_), .A2(new_n600_), .A3(new_n588_), .ZN(new_n612_));
  AOI21_X1  g0170(.A(new_n577_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g0171(.A1(new_n613_), .A2(new_n604_), .ZN(new_n614_));
  NAND3_X1  g0172(.A1(new_n607_), .A2(new_n603_), .A3(new_n614_), .ZN(new_n615_));
  OR2_X1    g0173(.A1(new_n507_), .A2(G214), .ZN(new_n616_));
  NAND2_X1  g0174(.A1(new_n616_), .A2(new_n509_), .ZN(new_n617_));
  INV_X1    g0175(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g0176(.A(G1480), .ZN(new_n619_));
  NOR2_X1   g0177(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g0178(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g0179(.A1(new_n618_), .A2(new_n619_), .ZN(new_n622_));
  NAND2_X1  g0180(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g0181(.A(G215), .ZN(new_n624_));
  AOI21_X1  g0182(.A(new_n573_), .B1(G18), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g0183(.A(G106), .ZN(new_n626_));
  NOR2_X1   g0184(.A1(new_n626_), .A2(KEYINPUT4), .ZN(new_n627_));
  OR2_X1    g0185(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g0186(.A1(new_n626_), .A2(KEYINPUT4), .ZN(new_n629_));
  OAI21_X1  g0187(.A(new_n625_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  AND2_X1   g0188(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g0189(.A1(new_n623_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g0190(.A(G209), .ZN(new_n633_));
  AOI21_X1  g0191(.A(new_n573_), .B1(G18), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g0192(.A(G1462), .ZN(new_n635_));
  NOR2_X1   g0193(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g0194(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g0195(.A1(new_n634_), .A2(new_n635_), .ZN(new_n638_));
  NAND2_X1  g0196(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g0197(.A(new_n509_), .B1(new_n507_), .B2(G216), .ZN(new_n640_));
  INV_X1    g0198(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g0199(.A(G1469), .ZN(new_n642_));
  NAND2_X1  g0200(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g0201(.A1(new_n640_), .A2(G1469), .ZN(new_n644_));
  NAND2_X1  g0202(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g0203(.A1(new_n639_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g0204(.A1(new_n632_), .A2(new_n646_), .ZN(new_n647_));
  OR2_X1    g0205(.A1(new_n507_), .A2(G213), .ZN(new_n648_));
  NAND2_X1  g0206(.A1(new_n648_), .A2(new_n509_), .ZN(new_n649_));
  INV_X1    g0207(.A(new_n649_), .ZN(new_n650_));
  INV_X1    g0208(.A(G1486), .ZN(new_n651_));
  NAND2_X1  g0209(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g0210(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g0211(.A1(new_n650_), .A2(new_n651_), .ZN(new_n654_));
  NOR2_X1   g0212(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g0213(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g0214(.A1(new_n647_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g0215(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g0216(.A1(G1492), .A2(G4528), .ZN(new_n659_));
  NOR2_X1   g0217(.A1(new_n659_), .A2(G38), .ZN(new_n660_));
  INV_X1    g0218(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g0219(.A(G38), .ZN(new_n662_));
  NAND3_X1  g0220(.A1(new_n662_), .A2(G1496), .A3(G4528), .ZN(new_n663_));
  NAND2_X1  g0221(.A1(G1496), .A2(G4528), .ZN(new_n664_));
  OAI21_X1  g0222(.A(G38), .B1(new_n659_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g0223(.A1(new_n661_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  NOR2_X1   g0224(.A1(new_n658_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g0225(.A1(new_n615_), .A2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g0226(.A(new_n668_), .B(KEYINPUT22), .Z(new_n669_));
  XNOR2_X1  g0227(.A(new_n665_), .B(KEYINPUT23), .ZN(new_n670_));
  NOR2_X1   g0228(.A1(new_n645_), .A2(new_n638_), .ZN(new_n671_));
  INV_X1    g0229(.A(new_n671_), .ZN(new_n672_));
  NAND2_X1  g0230(.A1(new_n643_), .A2(KEYINPUT24), .ZN(new_n673_));
  OR3_X1    g0231(.A1(new_n640_), .A2(KEYINPUT24), .A3(G1469), .ZN(new_n674_));
  NAND2_X1  g0232(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g0233(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g0234(.A(new_n631_), .B1(new_n672_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g0235(.A(new_n623_), .ZN(new_n678_));
  NAND3_X1  g0236(.A1(new_n677_), .A2(new_n655_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g0237(.A1(new_n625_), .A2(new_n626_), .ZN(new_n680_));
  AOI21_X1  g0238(.A(new_n620_), .B1(new_n622_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g0239(.A(new_n654_), .ZN(new_n682_));
  AOI21_X1  g0240(.A(new_n653_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g0241(.A1(new_n679_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g0242(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g0243(.A(new_n670_), .B1(new_n685_), .B2(new_n666_), .ZN(new_n686_));
  NOR2_X1   g0244(.A1(new_n669_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g0245(.A1(new_n507_), .A2(G103), .ZN(new_n688_));
  INV_X1    g0246(.A(G235), .ZN(new_n689_));
  OAI21_X1  g0247(.A(new_n688_), .B1(new_n507_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g0248(.A(new_n690_), .ZN(new_n691_));
  NOR2_X1   g0249(.A1(new_n691_), .A2(G3723), .ZN(new_n692_));
  NAND2_X1  g0250(.A1(new_n507_), .A2(G23), .ZN(new_n693_));
  INV_X1    g0251(.A(G236), .ZN(new_n694_));
  OAI21_X1  g0252(.A(new_n693_), .B1(new_n507_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g0253(.A(G3717), .ZN(new_n696_));
  NAND2_X1  g0254(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g0255(.A1(new_n507_), .A2(G26), .ZN(new_n698_));
  NAND2_X1  g0256(.A1(G18), .A2(G237), .ZN(new_n699_));
  NAND2_X1  g0257(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g0258(.A(G3711), .ZN(new_n701_));
  NAND2_X1  g0259(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g0260(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g0261(.A1(new_n698_), .A2(G3711), .A3(new_n699_), .ZN(new_n704_));
  NAND2_X1  g0262(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g0263(.A(KEYINPUT12), .ZN(new_n706_));
  NAND2_X1  g0264(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g0265(.A1(new_n700_), .A2(KEYINPUT12), .A3(G3711), .ZN(new_n708_));
  AND2_X1   g0266(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g0267(.A(KEYINPUT13), .B1(G18), .B2(G238), .ZN(new_n710_));
  NAND2_X1  g0268(.A1(new_n507_), .A2(G29), .ZN(new_n711_));
  NAND2_X1  g0269(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g0270(.A1(KEYINPUT13), .A2(G18), .A3(G238), .ZN(new_n713_));
  NAND2_X1  g0271(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g0272(.A(KEYINPUT14), .B(G3705), .ZN(new_n715_));
  NAND2_X1  g0273(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g0274(.A(G3705), .ZN(new_n717_));
  NAND3_X1  g0275(.A1(new_n712_), .A2(new_n717_), .A3(new_n713_), .ZN(new_n718_));
  NAND3_X1  g0276(.A1(new_n716_), .A2(new_n501_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g0277(.A1(new_n718_), .A2(KEYINPUT15), .ZN(new_n720_));
  INV_X1    g0278(.A(KEYINPUT15), .ZN(new_n721_));
  NAND4_X1  g0279(.A1(new_n712_), .A2(new_n721_), .A3(new_n717_), .A4(new_n713_), .ZN(new_n722_));
  NAND2_X1  g0280(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g0281(.A1(new_n719_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g0282(.A(new_n703_), .B1(new_n709_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g0283(.A(KEYINPUT11), .B(G3717), .ZN(new_n726_));
  NAND2_X1  g0284(.A1(new_n695_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g0285(.A(KEYINPUT11), .ZN(new_n728_));
  NOR2_X1   g0286(.A1(new_n728_), .A2(new_n696_), .ZN(new_n729_));
  OAI21_X1  g0287(.A(new_n727_), .B1(new_n695_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g0288(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g0289(.A(new_n697_), .B1(new_n725_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g0290(.A1(new_n691_), .A2(G3723), .ZN(new_n733_));
  AOI21_X1  g0291(.A(new_n692_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g0292(.A1(new_n707_), .A2(new_n708_), .A3(new_n730_), .ZN(new_n735_));
  INV_X1    g0293(.A(new_n692_), .ZN(new_n736_));
  NAND2_X1  g0294(.A1(new_n736_), .A2(new_n733_), .ZN(new_n737_));
  NAND3_X1  g0295(.A1(new_n716_), .A2(new_n504_), .A3(new_n718_), .ZN(new_n738_));
  NOR3_X1   g0296(.A1(new_n735_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g0297(.A1(new_n739_), .A2(G4526), .ZN(new_n740_));
  NAND2_X1  g0298(.A1(new_n734_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g0299(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g0300(.A1(new_n507_), .A2(G124), .ZN(new_n743_));
  NAND2_X1  g0301(.A1(G18), .A2(G232), .ZN(new_n744_));
  AND2_X1   g0302(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OR2_X1    g0303(.A1(new_n745_), .A2(G3743), .ZN(new_n746_));
  NAND2_X1  g0304(.A1(new_n745_), .A2(G3743), .ZN(new_n747_));
  NAND2_X1  g0305(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g0306(.A(new_n748_), .B(KEYINPUT16), .ZN(new_n749_));
  AND2_X1   g0307(.A1(new_n507_), .A2(G130), .ZN(new_n750_));
  AOI21_X1  g0308(.A(new_n750_), .B1(G18), .B2(G234), .ZN(new_n751_));
  NAND2_X1  g0309(.A1(new_n751_), .A2(G3729), .ZN(new_n752_));
  INV_X1    g0310(.A(new_n752_), .ZN(new_n753_));
  NOR2_X1   g0311(.A1(new_n751_), .A2(G3729), .ZN(new_n754_));
  NOR2_X1   g0312(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g0313(.A1(new_n507_), .A2(G127), .ZN(new_n756_));
  NAND2_X1  g0314(.A1(G18), .A2(G233), .ZN(new_n757_));
  AND2_X1   g0315(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OR2_X1    g0316(.A1(new_n758_), .A2(G3737), .ZN(new_n759_));
  NAND2_X1  g0317(.A1(new_n758_), .A2(G3737), .ZN(new_n760_));
  NAND2_X1  g0318(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g0319(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g0320(.A1(new_n507_), .A2(G100), .ZN(new_n763_));
  NAND2_X1  g0321(.A1(G18), .A2(G231), .ZN(new_n764_));
  AND2_X1   g0322(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OR2_X1    g0323(.A1(new_n765_), .A2(G3749), .ZN(new_n766_));
  NAND2_X1  g0324(.A1(new_n765_), .A2(G3749), .ZN(new_n767_));
  NAND4_X1  g0325(.A1(new_n755_), .A2(new_n762_), .A3(new_n766_), .A4(new_n767_), .ZN(new_n768_));
  NOR3_X1   g0326(.A1(new_n742_), .A2(new_n749_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g0327(.A(new_n759_), .ZN(new_n770_));
  NAND2_X1  g0328(.A1(new_n754_), .A2(new_n760_), .ZN(new_n771_));
  NOR3_X1   g0329(.A1(new_n749_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g0330(.A(KEYINPUT17), .ZN(new_n773_));
  XNOR2_X1  g0331(.A(new_n746_), .B(new_n773_), .ZN(new_n774_));
  OAI21_X1  g0332(.A(new_n774_), .B1(new_n748_), .B2(new_n759_), .ZN(new_n775_));
  OAI21_X1  g0333(.A(new_n767_), .B1(new_n772_), .B2(new_n775_), .ZN(new_n776_));
  AND2_X1   g0334(.A1(new_n776_), .A2(new_n766_), .ZN(new_n777_));
  INV_X1    g0335(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g0336(.A1(new_n769_), .A2(new_n778_), .ZN(new_n779_));
  MUX2_X1   g0337(.A(G47), .B(G223), .S(G18), .Z(new_n780_));
  INV_X1    g0338(.A(G4415), .ZN(new_n781_));
  OR2_X1    g0339(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g0340(.A1(new_n780_), .A2(new_n781_), .ZN(new_n783_));
  NAND2_X1  g0341(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g0342(.A(G118), .ZN(new_n785_));
  NOR2_X1   g0343(.A1(new_n785_), .A2(G18), .ZN(new_n786_));
  INV_X1    g0344(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g0345(.A(G217), .ZN(new_n788_));
  OAI21_X1  g0346(.A(new_n787_), .B1(new_n507_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g0347(.A(G4394), .ZN(new_n790_));
  NAND2_X1  g0348(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g0349(.A(new_n786_), .B1(G18), .B2(G217), .ZN(new_n792_));
  NAND2_X1  g0350(.A1(new_n792_), .A2(G4394), .ZN(new_n793_));
  NAND2_X1  g0351(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g0352(.A1(new_n507_), .A2(G97), .ZN(new_n795_));
  NAND2_X1  g0353(.A1(G18), .A2(G226), .ZN(new_n796_));
  NAND2_X1  g0354(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g0355(.A(G4400), .ZN(new_n798_));
  NAND2_X1  g0356(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g0357(.A1(new_n795_), .A2(G4400), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g0358(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g0359(.A1(new_n794_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g0360(.A1(new_n507_), .A2(G94), .ZN(new_n803_));
  NAND2_X1  g0361(.A1(G18), .A2(G225), .ZN(new_n804_));
  NAND2_X1  g0362(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g0363(.A(new_n805_), .ZN(new_n806_));
  INV_X1    g0364(.A(G4405), .ZN(new_n807_));
  NAND2_X1  g0365(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g0366(.A1(new_n805_), .A2(G4405), .ZN(new_n809_));
  NAND2_X1  g0367(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g0368(.A1(new_n507_), .A2(G121), .ZN(new_n811_));
  INV_X1    g0369(.A(G224), .ZN(new_n812_));
  OAI21_X1  g0370(.A(new_n811_), .B1(new_n507_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g0371(.A(new_n813_), .B(G4410), .ZN(new_n814_));
  NAND3_X1  g0372(.A1(new_n802_), .A2(new_n810_), .A3(new_n814_), .ZN(new_n815_));
  NOR3_X1   g0373(.A1(new_n779_), .A2(new_n784_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g0374(.A1(new_n507_), .A2(G32), .ZN(new_n817_));
  NAND2_X1  g0375(.A1(G18), .A2(G221), .ZN(new_n818_));
  NAND2_X1  g0376(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g0377(.A(G4427), .ZN(new_n820_));
  NAND2_X1  g0378(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g0379(.A1(new_n817_), .A2(G4427), .A3(new_n818_), .ZN(new_n822_));
  AND2_X1   g0380(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g0381(.A(new_n823_), .B(KEYINPUT18), .ZN(new_n824_));
  INV_X1    g0382(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g0383(.A1(new_n507_), .A2(G50), .ZN(new_n826_));
  NAND2_X1  g0384(.A1(G18), .A2(G220), .ZN(new_n827_));
  AND2_X1   g0385(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OR2_X1    g0386(.A1(new_n828_), .A2(G4432), .ZN(new_n829_));
  NAND2_X1  g0387(.A1(new_n828_), .A2(G4432), .ZN(new_n830_));
  AND2_X1   g0388(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g0389(.A(KEYINPUT19), .B(G4420), .ZN(new_n832_));
  NAND2_X1  g0390(.A1(new_n507_), .A2(G35), .ZN(new_n833_));
  NAND2_X1  g0391(.A1(G18), .A2(G222), .ZN(new_n834_));
  NAND2_X1  g0392(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g0393(.A(new_n832_), .B(new_n835_), .ZN(new_n836_));
  NAND2_X1  g0394(.A1(new_n507_), .A2(G66), .ZN(new_n837_));
  INV_X1    g0395(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g0396(.A(new_n838_), .B1(G18), .B2(G219), .ZN(new_n839_));
  OR2_X1    g0397(.A1(new_n839_), .A2(G4437), .ZN(new_n840_));
  NAND2_X1  g0398(.A1(new_n839_), .A2(G4437), .ZN(new_n841_));
  NAND4_X1  g0399(.A1(new_n831_), .A2(new_n836_), .A3(new_n840_), .A4(new_n841_), .ZN(new_n842_));
  NOR2_X1   g0400(.A1(new_n825_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g0401(.A1(new_n816_), .A2(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g0402(.A(new_n799_), .B(KEYINPUT26), .ZN(new_n845_));
  NAND3_X1  g0403(.A1(new_n845_), .A2(new_n810_), .A3(new_n814_), .ZN(new_n846_));
  INV_X1    g0404(.A(KEYINPUT27), .ZN(new_n847_));
  OR2_X1    g0405(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g0406(.A1(new_n806_), .A2(G4405), .ZN(new_n849_));
  INV_X1    g0407(.A(new_n849_), .ZN(new_n850_));
  INV_X1    g0408(.A(new_n801_), .ZN(new_n851_));
  NOR2_X1   g0409(.A1(new_n792_), .A2(G4394), .ZN(new_n852_));
  NAND2_X1  g0410(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g0411(.A(new_n810_), .ZN(new_n854_));
  OAI21_X1  g0412(.A(new_n850_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g0413(.A1(new_n855_), .A2(new_n814_), .ZN(new_n856_));
  AOI21_X1  g0414(.A(new_n784_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g0415(.A(new_n847_), .B1(new_n846_), .B2(new_n784_), .ZN(new_n858_));
  XOR2_X1   g0416(.A(new_n783_), .B(KEYINPUT25), .Z(new_n859_));
  INV_X1    g0417(.A(G4410), .ZN(new_n860_));
  NAND2_X1  g0418(.A1(new_n813_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g0419(.A(new_n784_), .B(KEYINPUT28), .ZN(new_n862_));
  OAI211_X1 g0420(.A(new_n858_), .B(new_n859_), .C1(new_n861_), .C2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g0421(.A1(new_n857_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g0422(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g0423(.A1(new_n865_), .A2(new_n843_), .ZN(new_n866_));
  XNOR2_X1  g0424(.A(new_n866_), .B(KEYINPUT29), .ZN(new_n867_));
  XOR2_X1   g0425(.A(new_n821_), .B(KEYINPUT30), .Z(new_n868_));
  NAND2_X1  g0426(.A1(new_n868_), .A2(new_n829_), .ZN(new_n869_));
  NAND2_X1  g0427(.A1(new_n869_), .A2(new_n830_), .ZN(new_n870_));
  INV_X1    g0428(.A(new_n835_), .ZN(new_n871_));
  NOR2_X1   g0429(.A1(new_n871_), .A2(G4420), .ZN(new_n872_));
  NAND3_X1  g0430(.A1(new_n831_), .A2(new_n823_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g0431(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g0432(.A1(new_n874_), .A2(new_n841_), .ZN(new_n875_));
  NAND2_X1  g0433(.A1(new_n875_), .A2(new_n840_), .ZN(new_n876_));
  NOR2_X1   g0434(.A1(new_n867_), .A2(new_n876_), .ZN(new_n877_));
  AND2_X1   g0435(.A1(new_n844_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g0436(.A(new_n566_), .ZN(new_n879_));
  NAND2_X1  g0437(.A1(new_n526_), .A2(new_n530_), .ZN(new_n880_));
  AND2_X1   g0438(.A1(new_n555_), .A2(new_n558_), .ZN(new_n881_));
  INV_X1    g0439(.A(new_n552_), .ZN(new_n882_));
  AOI21_X1  g0440(.A(KEYINPUT8), .B1(new_n556_), .B2(new_n547_), .ZN(new_n883_));
  OAI21_X1  g0441(.A(G2230), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g0442(.A(new_n880_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g0443(.A(G2211), .ZN(new_n886_));
  INV_X1    g0444(.A(new_n539_), .ZN(new_n887_));
  AOI211_X1 g0445(.A(new_n886_), .B(new_n887_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n888_));
  NAND2_X1  g0446(.A1(new_n519_), .A2(new_n532_), .ZN(new_n889_));
  NOR3_X1   g0447(.A1(new_n888_), .A2(new_n540_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g0448(.A1(new_n885_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g0449(.A1(new_n879_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g0450(.A1(new_n606_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g0451(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g0452(.A1(new_n894_), .A2(new_n667_), .ZN(new_n895_));
  OAI21_X1  g0453(.A(new_n687_), .B1(new_n878_), .B2(new_n895_), .ZN(G246));
  OAI21_X1  g0454(.A(new_n509_), .B1(new_n507_), .B2(G173), .ZN(new_n897_));
  XNOR2_X1  g0455(.A(new_n897_), .B(KEYINPUT38), .ZN(new_n898_));
  INV_X1    g0456(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g0457(.A1(new_n507_), .A2(G2256), .ZN(new_n900_));
  AOI21_X1  g0458(.A(new_n900_), .B1(new_n507_), .B2(G110), .ZN(new_n901_));
  OR2_X1    g0459(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g0460(.A(new_n902_), .B(KEYINPUT47), .ZN(new_n903_));
  OAI21_X1  g0461(.A(new_n509_), .B1(new_n507_), .B2(G174), .ZN(new_n904_));
  NAND2_X1  g0462(.A1(new_n507_), .A2(G109), .ZN(new_n905_));
  NAND2_X1  g0463(.A1(new_n576_), .A2(G18), .ZN(new_n906_));
  AND2_X1   g0464(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  AOI22_X1  g0465(.A1(new_n899_), .A2(new_n901_), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g0466(.A1(new_n902_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g0467(.A1(new_n907_), .A2(new_n904_), .ZN(new_n910_));
  OR2_X1    g0468(.A1(new_n507_), .A2(G175), .ZN(new_n911_));
  NAND2_X1  g0469(.A1(new_n911_), .A2(new_n509_), .ZN(new_n912_));
  INV_X1    g0470(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g0471(.A1(new_n507_), .A2(G86), .ZN(new_n914_));
  OAI21_X1  g0472(.A(new_n914_), .B1(new_n507_), .B2(G2247), .ZN(new_n915_));
  AOI21_X1  g0473(.A(new_n910_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g0474(.A(new_n916_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n917_));
  OR2_X1    g0475(.A1(new_n909_), .A2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g0476(.A(new_n509_), .B1(new_n507_), .B2(G176), .ZN(new_n919_));
  INV_X1    g0477(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g0478(.A1(new_n507_), .A2(G63), .ZN(new_n921_));
  OAI21_X1  g0479(.A(new_n921_), .B1(new_n507_), .B2(G2239), .ZN(new_n922_));
  NAND2_X1  g0480(.A1(new_n920_), .A2(new_n922_), .ZN(new_n923_));
  OAI221_X1 g0481(.A(new_n903_), .B1(new_n909_), .B2(new_n916_), .C1(new_n918_), .C2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g0482(.A1(new_n507_), .A2(G64), .ZN(new_n925_));
  OAI21_X1  g0483(.A(new_n925_), .B1(new_n507_), .B2(G2236), .ZN(new_n926_));
  OAI21_X1  g0484(.A(new_n509_), .B1(new_n507_), .B2(G177), .ZN(new_n927_));
  XNOR2_X1  g0485(.A(new_n926_), .B(new_n927_), .ZN(new_n928_));
  INV_X1    g0486(.A(G178), .ZN(new_n929_));
  OAI21_X1  g0487(.A(new_n556_), .B1(new_n507_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g0488(.A1(new_n507_), .A2(G85), .ZN(new_n931_));
  OAI21_X1  g0489(.A(new_n931_), .B1(new_n507_), .B2(G2230), .ZN(new_n932_));
  AND3_X1   g0490(.A1(new_n928_), .A2(new_n930_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g0491(.A(KEYINPUT37), .ZN(new_n934_));
  INV_X1    g0492(.A(new_n522_), .ZN(new_n935_));
  AOI21_X1  g0493(.A(new_n935_), .B1(G18), .B2(G179), .ZN(new_n936_));
  INV_X1    g0494(.A(new_n936_), .ZN(new_n937_));
  NAND2_X1  g0495(.A1(new_n507_), .A2(G84), .ZN(new_n938_));
  NAND2_X1  g0496(.A1(new_n525_), .A2(G18), .ZN(new_n939_));
  AND2_X1   g0497(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g0498(.A(new_n940_), .ZN(new_n941_));
  OAI22_X1  g0499(.A1(new_n928_), .A2(new_n934_), .B1(new_n937_), .B2(new_n941_), .ZN(new_n942_));
  AOI21_X1  g0500(.A(new_n942_), .B1(new_n934_), .B2(new_n928_), .ZN(new_n943_));
  XOR2_X1   g0501(.A(new_n930_), .B(new_n932_), .Z(new_n944_));
  INV_X1    g0502(.A(new_n944_), .ZN(new_n945_));
  NOR2_X1   g0503(.A1(new_n516_), .A2(G18), .ZN(new_n946_));
  AOI21_X1  g0504(.A(new_n946_), .B1(G18), .B2(G180), .ZN(new_n947_));
  INV_X1    g0505(.A(new_n947_), .ZN(new_n948_));
  NAND2_X1  g0506(.A1(new_n507_), .A2(G83), .ZN(new_n949_));
  OAI21_X1  g0507(.A(new_n949_), .B1(new_n507_), .B2(G2218), .ZN(new_n950_));
  AOI22_X1  g0508(.A1(new_n937_), .A2(new_n941_), .B1(new_n948_), .B2(new_n950_), .ZN(new_n951_));
  NOR2_X1   g0509(.A1(new_n945_), .A2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g0510(.A1(new_n943_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g0511(.A(new_n926_), .ZN(new_n954_));
  OAI21_X1  g0512(.A(new_n953_), .B1(new_n927_), .B2(new_n954_), .ZN(new_n955_));
  OR2_X1    g0513(.A1(new_n948_), .A2(new_n950_), .ZN(new_n956_));
  AND3_X1   g0514(.A1(new_n943_), .A2(new_n956_), .A3(new_n951_), .ZN(new_n957_));
  NAND2_X1  g0515(.A1(new_n507_), .A2(G65), .ZN(new_n958_));
  OAI21_X1  g0516(.A(new_n958_), .B1(new_n507_), .B2(G2211), .ZN(new_n959_));
  XOR2_X1   g0517(.A(new_n959_), .B(KEYINPUT36), .Z(new_n960_));
  AOI22_X1  g0518(.A1(new_n535_), .A2(new_n537_), .B1(G18), .B2(G171), .ZN(new_n961_));
  INV_X1    g0519(.A(new_n961_), .ZN(new_n962_));
  NAND2_X1  g0520(.A1(new_n960_), .A2(new_n962_), .ZN(new_n963_));
  NOR2_X1   g0521(.A1(new_n963_), .A2(new_n945_), .ZN(new_n964_));
  XOR2_X1   g0522(.A(new_n964_), .B(KEYINPUT45), .Z(new_n965_));
  AOI21_X1  g0523(.A(new_n955_), .B1(new_n957_), .B2(new_n965_), .ZN(new_n966_));
  INV_X1    g0524(.A(KEYINPUT46), .ZN(new_n967_));
  AOI21_X1  g0525(.A(new_n933_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g0526(.A(new_n968_), .B1(new_n967_), .B2(new_n966_), .ZN(new_n969_));
  XNOR2_X1  g0527(.A(new_n920_), .B(new_n922_), .ZN(new_n970_));
  NOR2_X1   g0528(.A1(new_n918_), .A2(new_n970_), .ZN(new_n971_));
  AOI21_X1  g0529(.A(new_n924_), .B1(new_n969_), .B2(new_n971_), .ZN(new_n972_));
  NAND2_X1  g0530(.A1(new_n507_), .A2(G112), .ZN(new_n973_));
  OAI21_X1  g0531(.A(new_n973_), .B1(new_n507_), .B2(G1480), .ZN(new_n974_));
  XOR2_X1   g0532(.A(new_n974_), .B(KEYINPUT34), .Z(new_n975_));
  OR2_X1    g0533(.A1(new_n507_), .A2(G167), .ZN(new_n976_));
  NAND2_X1  g0534(.A1(new_n976_), .A2(new_n509_), .ZN(new_n977_));
  NOR2_X1   g0535(.A1(new_n975_), .A2(new_n977_), .ZN(new_n978_));
  OAI21_X1  g0536(.A(new_n509_), .B1(new_n507_), .B2(G166), .ZN(new_n979_));
  INV_X1    g0537(.A(new_n979_), .ZN(new_n980_));
  NOR2_X1   g0538(.A1(new_n507_), .A2(G1486), .ZN(new_n981_));
  AOI21_X1  g0539(.A(new_n981_), .B1(new_n507_), .B2(G88), .ZN(new_n982_));
  INV_X1    g0540(.A(new_n982_), .ZN(new_n983_));
  AOI21_X1  g0541(.A(new_n978_), .B1(new_n980_), .B2(new_n983_), .ZN(new_n984_));
  NOR2_X1   g0542(.A1(new_n983_), .A2(new_n980_), .ZN(new_n985_));
  INV_X1    g0543(.A(new_n985_), .ZN(new_n986_));
  NAND2_X1  g0544(.A1(new_n975_), .A2(new_n977_), .ZN(new_n987_));
  NAND3_X1  g0545(.A1(new_n984_), .A2(new_n986_), .A3(new_n987_), .ZN(new_n988_));
  NAND2_X1  g0546(.A1(new_n507_), .A2(G87), .ZN(new_n989_));
  OAI21_X1  g0547(.A(new_n989_), .B1(new_n507_), .B2(G106), .ZN(new_n990_));
  OAI21_X1  g0548(.A(new_n509_), .B1(new_n507_), .B2(G168), .ZN(new_n991_));
  XNOR2_X1  g0549(.A(new_n990_), .B(new_n991_), .ZN(new_n992_));
  NAND2_X1  g0550(.A1(new_n507_), .A2(G111), .ZN(new_n993_));
  OAI21_X1  g0551(.A(new_n993_), .B1(new_n507_), .B2(G1469), .ZN(new_n994_));
  OR2_X1    g0552(.A1(new_n507_), .A2(G169), .ZN(new_n995_));
  NAND3_X1  g0553(.A1(new_n994_), .A2(new_n509_), .A3(new_n995_), .ZN(new_n996_));
  INV_X1    g0554(.A(new_n994_), .ZN(new_n997_));
  NAND2_X1  g0555(.A1(new_n995_), .A2(new_n509_), .ZN(new_n998_));
  NAND2_X1  g0556(.A1(new_n997_), .A2(new_n998_), .ZN(new_n999_));
  NAND3_X1  g0557(.A1(new_n992_), .A2(new_n996_), .A3(new_n999_), .ZN(new_n1000_));
  NAND2_X1  g0558(.A1(new_n507_), .A2(G113), .ZN(new_n1001_));
  OAI21_X1  g0559(.A(new_n1001_), .B1(new_n507_), .B2(G1462), .ZN(new_n1002_));
  XNOR2_X1  g0560(.A(new_n1002_), .B(new_n509_), .ZN(new_n1003_));
  NOR3_X1   g0561(.A1(new_n988_), .A2(new_n1000_), .A3(new_n1003_), .ZN(new_n1004_));
  INV_X1    g0562(.A(G1455), .ZN(new_n1005_));
  NAND2_X1  g0563(.A1(new_n1005_), .A2(G4528), .ZN(new_n1006_));
  XNOR2_X1  g0564(.A(new_n1006_), .B(KEYINPUT35), .ZN(new_n1007_));
  INV_X1    g0565(.A(G4528), .ZN(new_n1008_));
  NOR3_X1   g0566(.A1(new_n1007_), .A2(G2204), .A3(new_n1008_), .ZN(new_n1009_));
  INV_X1    g0567(.A(G2204), .ZN(new_n1010_));
  AOI21_X1  g0568(.A(G38), .B1(new_n1010_), .B2(G4528), .ZN(new_n1011_));
  AOI22_X1  g0569(.A1(new_n1009_), .A2(G38), .B1(new_n1007_), .B2(new_n1011_), .ZN(new_n1012_));
  INV_X1    g0570(.A(new_n1012_), .ZN(new_n1013_));
  NAND2_X1  g0571(.A1(new_n1004_), .A2(new_n1013_), .ZN(new_n1014_));
  NOR2_X1   g0572(.A1(new_n972_), .A2(new_n1014_), .ZN(new_n1015_));
  XNOR2_X1  g0573(.A(new_n1015_), .B(KEYINPUT48), .ZN(new_n1016_));
  INV_X1    g0574(.A(G190), .ZN(new_n1017_));
  OAI21_X1  g0575(.A(new_n826_), .B1(new_n507_), .B2(new_n1017_), .ZN(new_n1018_));
  NAND2_X1  g0576(.A1(new_n507_), .A2(G61), .ZN(new_n1019_));
  OAI21_X1  g0577(.A(new_n1019_), .B1(new_n507_), .B2(G4432), .ZN(new_n1020_));
  NAND2_X1  g0578(.A1(new_n1018_), .A2(new_n1020_), .ZN(new_n1021_));
  INV_X1    g0579(.A(G191), .ZN(new_n1022_));
  OAI21_X1  g0580(.A(new_n817_), .B1(new_n507_), .B2(new_n1022_), .ZN(new_n1023_));
  XNOR2_X1  g0581(.A(new_n1023_), .B(KEYINPUT43), .ZN(new_n1024_));
  NAND2_X1  g0582(.A1(new_n507_), .A2(G60), .ZN(new_n1025_));
  OAI21_X1  g0583(.A(new_n1025_), .B1(new_n507_), .B2(G4427), .ZN(new_n1026_));
  NAND2_X1  g0584(.A1(new_n1024_), .A2(new_n1026_), .ZN(new_n1027_));
  NOR2_X1   g0585(.A1(new_n1024_), .A2(new_n1026_), .ZN(new_n1028_));
  INV_X1    g0586(.A(new_n833_), .ZN(new_n1029_));
  AOI21_X1  g0587(.A(new_n1029_), .B1(G18), .B2(G192), .ZN(new_n1030_));
  NOR2_X1   g0588(.A1(new_n507_), .A2(G4420), .ZN(new_n1031_));
  AOI21_X1  g0589(.A(new_n1031_), .B1(new_n507_), .B2(G79), .ZN(new_n1032_));
  OR2_X1    g0590(.A1(new_n1030_), .A2(new_n1032_), .ZN(new_n1033_));
  OAI211_X1 g0591(.A(new_n1021_), .B(new_n1027_), .C1(new_n1028_), .C2(new_n1033_), .ZN(new_n1034_));
  OR2_X1    g0592(.A1(new_n1018_), .A2(new_n1020_), .ZN(new_n1035_));
  NAND2_X1  g0593(.A1(new_n507_), .A2(G62), .ZN(new_n1036_));
  OAI21_X1  g0594(.A(new_n1036_), .B1(new_n507_), .B2(G4437), .ZN(new_n1037_));
  XOR2_X1   g0595(.A(new_n1037_), .B(KEYINPUT42), .Z(new_n1038_));
  AOI21_X1  g0596(.A(new_n838_), .B1(G18), .B2(G189), .ZN(new_n1039_));
  NAND2_X1  g0597(.A1(new_n1038_), .A2(new_n1039_), .ZN(new_n1040_));
  NAND3_X1  g0598(.A1(new_n1034_), .A2(new_n1035_), .A3(new_n1040_), .ZN(new_n1041_));
  OR2_X1    g0599(.A1(new_n1038_), .A2(new_n1039_), .ZN(new_n1042_));
  NAND2_X1  g0600(.A1(new_n1041_), .A2(new_n1042_), .ZN(new_n1043_));
  NAND3_X1  g0601(.A1(new_n1042_), .A2(new_n1027_), .A3(new_n1040_), .ZN(new_n1044_));
  NAND2_X1  g0602(.A1(new_n1030_), .A2(new_n1032_), .ZN(new_n1045_));
  NAND4_X1  g0603(.A1(new_n1033_), .A2(new_n1021_), .A3(new_n1035_), .A4(new_n1045_), .ZN(new_n1046_));
  NOR3_X1   g0604(.A1(new_n1044_), .A2(new_n1028_), .A3(new_n1046_), .ZN(new_n1047_));
  XOR2_X1   g0605(.A(new_n1047_), .B(KEYINPUT44), .Z(new_n1048_));
  NAND2_X1  g0606(.A1(new_n507_), .A2(G80), .ZN(new_n1049_));
  OAI21_X1  g0607(.A(new_n1049_), .B1(new_n507_), .B2(G4415), .ZN(new_n1050_));
  INV_X1    g0608(.A(new_n1050_), .ZN(new_n1051_));
  AND2_X1   g0609(.A1(G18), .A2(G193), .ZN(new_n1052_));
  AOI21_X1  g0610(.A(new_n1052_), .B1(new_n507_), .B2(G47), .ZN(new_n1053_));
  NOR2_X1   g0611(.A1(new_n1051_), .A2(new_n1053_), .ZN(new_n1054_));
  INV_X1    g0612(.A(G194), .ZN(new_n1055_));
  OAI21_X1  g0613(.A(new_n811_), .B1(new_n507_), .B2(new_n1055_), .ZN(new_n1056_));
  XNOR2_X1  g0614(.A(new_n1056_), .B(KEYINPUT40), .ZN(new_n1057_));
  OR3_X1    g0615(.A1(new_n507_), .A2(KEYINPUT39), .A3(G4410), .ZN(new_n1058_));
  NAND2_X1  g0616(.A1(new_n507_), .A2(G81), .ZN(new_n1059_));
  OAI21_X1  g0617(.A(KEYINPUT39), .B1(new_n507_), .B2(G4410), .ZN(new_n1060_));
  NAND3_X1  g0618(.A1(new_n1058_), .A2(new_n1059_), .A3(new_n1060_), .ZN(new_n1061_));
  NAND2_X1  g0619(.A1(new_n1057_), .A2(new_n1061_), .ZN(new_n1062_));
  INV_X1    g0620(.A(G195), .ZN(new_n1063_));
  OAI21_X1  g0621(.A(new_n803_), .B1(new_n507_), .B2(new_n1063_), .ZN(new_n1064_));
  NAND2_X1  g0622(.A1(new_n507_), .A2(G59), .ZN(new_n1065_));
  OAI21_X1  g0623(.A(new_n1065_), .B1(new_n507_), .B2(G4405), .ZN(new_n1066_));
  NAND2_X1  g0624(.A1(new_n1064_), .A2(new_n1066_), .ZN(new_n1067_));
  NAND2_X1  g0625(.A1(new_n798_), .A2(G18), .ZN(new_n1068_));
  AOI22_X1  g0626(.A1(new_n1068_), .A2(KEYINPUT41), .B1(new_n507_), .B2(G78), .ZN(new_n1069_));
  OAI21_X1  g0627(.A(new_n1069_), .B1(KEYINPUT41), .B2(new_n1068_), .ZN(new_n1070_));
  INV_X1    g0628(.A(G196), .ZN(new_n1071_));
  OAI21_X1  g0629(.A(new_n795_), .B1(new_n507_), .B2(new_n1071_), .ZN(new_n1072_));
  INV_X1    g0630(.A(G187), .ZN(new_n1073_));
  OAI21_X1  g0631(.A(new_n787_), .B1(new_n507_), .B2(new_n1073_), .ZN(new_n1074_));
  NAND2_X1  g0632(.A1(new_n507_), .A2(G77), .ZN(new_n1075_));
  OAI21_X1  g0633(.A(new_n1075_), .B1(new_n507_), .B2(G4394), .ZN(new_n1076_));
  AOI22_X1  g0634(.A1(new_n1070_), .A2(new_n1072_), .B1(new_n1074_), .B2(new_n1076_), .ZN(new_n1077_));
  OAI22_X1  g0635(.A1(new_n1070_), .A2(new_n1072_), .B1(new_n1064_), .B2(new_n1066_), .ZN(new_n1078_));
  OAI211_X1 g0636(.A(new_n1062_), .B(new_n1067_), .C1(new_n1077_), .C2(new_n1078_), .ZN(new_n1079_));
  OR2_X1    g0637(.A1(new_n1057_), .A2(new_n1061_), .ZN(new_n1080_));
  NAND2_X1  g0638(.A1(new_n1051_), .A2(new_n1053_), .ZN(new_n1081_));
  NAND3_X1  g0639(.A1(new_n1079_), .A2(new_n1080_), .A3(new_n1081_), .ZN(new_n1082_));
  NAND2_X1  g0640(.A1(new_n1082_), .A2(KEYINPUT51), .ZN(new_n1083_));
  NOR2_X1   g0641(.A1(new_n1067_), .A2(KEYINPUT51), .ZN(new_n1084_));
  NAND4_X1  g0642(.A1(new_n1080_), .A2(new_n1062_), .A3(new_n1081_), .A4(new_n1084_), .ZN(new_n1085_));
  AOI21_X1  g0643(.A(new_n1054_), .B1(new_n1083_), .B2(new_n1085_), .ZN(new_n1086_));
  INV_X1    g0644(.A(new_n1086_), .ZN(new_n1087_));
  AOI21_X1  g0645(.A(new_n1043_), .B1(new_n1048_), .B2(new_n1087_), .ZN(new_n1088_));
  OR2_X1    g0646(.A1(new_n960_), .A2(new_n962_), .ZN(new_n1089_));
  AND3_X1   g0647(.A1(new_n1089_), .A2(new_n963_), .A3(new_n944_), .ZN(new_n1090_));
  NAND3_X1  g0648(.A1(new_n971_), .A2(new_n957_), .A3(new_n1090_), .ZN(new_n1091_));
  OR2_X1    g0649(.A1(new_n1014_), .A2(new_n1091_), .ZN(new_n1092_));
  NOR2_X1   g0650(.A1(new_n1088_), .A2(new_n1092_), .ZN(new_n1093_));
  XOR2_X1   g0651(.A(new_n1093_), .B(KEYINPUT52), .Z(new_n1094_));
  INV_X1    g0652(.A(G200), .ZN(new_n1095_));
  OAI21_X1  g0653(.A(new_n763_), .B1(new_n507_), .B2(new_n1095_), .ZN(new_n1096_));
  NAND2_X1  g0654(.A1(new_n507_), .A2(G56), .ZN(new_n1097_));
  OAI21_X1  g0655(.A(new_n1097_), .B1(new_n507_), .B2(G3749), .ZN(new_n1098_));
  OAI211_X1 g0656(.A(new_n1081_), .B(new_n1067_), .C1(new_n1096_), .C2(new_n1098_), .ZN(new_n1099_));
  NOR2_X1   g0657(.A1(new_n1074_), .A2(new_n1076_), .ZN(new_n1100_));
  NOR3_X1   g0658(.A1(new_n1099_), .A2(new_n1054_), .A3(new_n1100_), .ZN(new_n1101_));
  NAND2_X1  g0659(.A1(new_n1101_), .A2(new_n1077_), .ZN(new_n1102_));
  NAND2_X1  g0660(.A1(new_n1080_), .A2(new_n1062_), .ZN(new_n1103_));
  NOR3_X1   g0661(.A1(new_n1102_), .A2(new_n1078_), .A3(new_n1103_), .ZN(new_n1104_));
  INV_X1    g0662(.A(G201), .ZN(new_n1105_));
  OAI21_X1  g0663(.A(new_n743_), .B1(new_n507_), .B2(new_n1105_), .ZN(new_n1106_));
  NAND2_X1  g0664(.A1(new_n507_), .A2(G55), .ZN(new_n1107_));
  OAI21_X1  g0665(.A(new_n1107_), .B1(new_n507_), .B2(G3743), .ZN(new_n1108_));
  NOR2_X1   g0666(.A1(new_n1106_), .A2(new_n1108_), .ZN(new_n1109_));
  INV_X1    g0667(.A(G202), .ZN(new_n1110_));
  OAI21_X1  g0668(.A(new_n756_), .B1(new_n507_), .B2(new_n1110_), .ZN(new_n1111_));
  NAND2_X1  g0669(.A1(new_n507_), .A2(G54), .ZN(new_n1112_));
  OAI21_X1  g0670(.A(new_n1112_), .B1(new_n507_), .B2(G3737), .ZN(new_n1113_));
  AOI21_X1  g0671(.A(new_n1109_), .B1(new_n1111_), .B2(new_n1113_), .ZN(new_n1114_));
  OAI21_X1  g0672(.A(new_n1114_), .B1(new_n1111_), .B2(new_n1113_), .ZN(new_n1115_));
  INV_X1    g0673(.A(G204), .ZN(new_n1116_));
  OAI21_X1  g0674(.A(new_n688_), .B1(new_n507_), .B2(new_n1116_), .ZN(new_n1117_));
  NAND2_X1  g0675(.A1(new_n507_), .A2(G73), .ZN(new_n1118_));
  OAI21_X1  g0676(.A(new_n1118_), .B1(new_n507_), .B2(G3723), .ZN(new_n1119_));
  NAND2_X1  g0677(.A1(new_n1117_), .A2(new_n1119_), .ZN(new_n1120_));
  MUX2_X1   g0678(.A(G130), .B(G203), .S(G18), .Z(new_n1121_));
  XNOR2_X1  g0679(.A(new_n1121_), .B(KEYINPUT31), .ZN(new_n1122_));
  OR2_X1    g0680(.A1(new_n507_), .A2(G3729), .ZN(new_n1123_));
  INV_X1    g0681(.A(G53), .ZN(new_n1124_));
  OAI21_X1  g0682(.A(new_n1123_), .B1(G18), .B2(new_n1124_), .ZN(new_n1125_));
  INV_X1    g0683(.A(new_n1125_), .ZN(new_n1126_));
  OAI21_X1  g0684(.A(new_n1120_), .B1(new_n1122_), .B2(new_n1126_), .ZN(new_n1127_));
  INV_X1    g0685(.A(G205), .ZN(new_n1128_));
  OAI21_X1  g0686(.A(new_n693_), .B1(new_n507_), .B2(new_n1128_), .ZN(new_n1129_));
  XNOR2_X1  g0687(.A(new_n1129_), .B(KEYINPUT32), .ZN(new_n1130_));
  NAND2_X1  g0688(.A1(new_n507_), .A2(G75), .ZN(new_n1131_));
  OAI21_X1  g0689(.A(new_n1131_), .B1(new_n507_), .B2(G3717), .ZN(new_n1132_));
  NAND2_X1  g0690(.A1(new_n1130_), .A2(new_n1132_), .ZN(new_n1133_));
  INV_X1    g0691(.A(G206), .ZN(new_n1134_));
  OAI21_X1  g0692(.A(new_n698_), .B1(new_n507_), .B2(new_n1134_), .ZN(new_n1135_));
  NAND2_X1  g0693(.A1(new_n507_), .A2(G76), .ZN(new_n1136_));
  OAI21_X1  g0694(.A(new_n1136_), .B1(new_n507_), .B2(G3711), .ZN(new_n1137_));
  INV_X1    g0695(.A(G207), .ZN(new_n1138_));
  OAI21_X1  g0696(.A(new_n711_), .B1(new_n507_), .B2(new_n1138_), .ZN(new_n1139_));
  NAND2_X1  g0697(.A1(new_n507_), .A2(G74), .ZN(new_n1140_));
  OAI21_X1  g0698(.A(new_n1140_), .B1(new_n507_), .B2(G3705), .ZN(new_n1141_));
  AOI22_X1  g0699(.A1(new_n1135_), .A2(new_n1137_), .B1(new_n1139_), .B2(new_n1141_), .ZN(new_n1142_));
  OR3_X1    g0700(.A1(G18), .A2(G41), .A3(G70), .ZN(new_n1143_));
  NAND3_X1  g0701(.A1(new_n507_), .A2(G41), .A3(G70), .ZN(new_n1144_));
  NAND4_X1  g0702(.A1(new_n1142_), .A2(G89), .A3(new_n1143_), .A4(new_n1144_), .ZN(new_n1145_));
  OR2_X1    g0703(.A1(new_n1135_), .A2(new_n1137_), .ZN(new_n1146_));
  OAI211_X1 g0704(.A(new_n1146_), .B(new_n1120_), .C1(new_n1139_), .C2(new_n1141_), .ZN(new_n1147_));
  OAI21_X1  g0705(.A(new_n1133_), .B1(new_n1145_), .B2(new_n1147_), .ZN(new_n1148_));
  NOR2_X1   g0706(.A1(new_n1117_), .A2(new_n1119_), .ZN(new_n1149_));
  INV_X1    g0707(.A(new_n1149_), .ZN(new_n1150_));
  NAND2_X1  g0708(.A1(new_n1148_), .A2(new_n1150_), .ZN(new_n1151_));
  NOR2_X1   g0709(.A1(new_n1139_), .A2(new_n1141_), .ZN(new_n1152_));
  OAI21_X1  g0710(.A(new_n1142_), .B1(new_n1152_), .B2(new_n1144_), .ZN(new_n1153_));
  OAI211_X1 g0711(.A(new_n1153_), .B(new_n1146_), .C1(KEYINPUT33), .C2(new_n1149_), .ZN(new_n1154_));
  INV_X1    g0712(.A(KEYINPUT33), .ZN(new_n1155_));
  AOI21_X1  g0713(.A(new_n1150_), .B1(new_n1133_), .B2(new_n1155_), .ZN(new_n1156_));
  OAI21_X1  g0714(.A(new_n1151_), .B1(new_n1154_), .B2(new_n1156_), .ZN(new_n1157_));
  OR2_X1    g0715(.A1(new_n1130_), .A2(new_n1132_), .ZN(new_n1158_));
  AOI21_X1  g0716(.A(new_n1127_), .B1(new_n1157_), .B2(new_n1158_), .ZN(new_n1159_));
  AOI211_X1 g0717(.A(new_n1115_), .B(new_n1159_), .C1(new_n1122_), .C2(new_n1126_), .ZN(new_n1160_));
  NAND2_X1  g0718(.A1(new_n1106_), .A2(new_n1108_), .ZN(new_n1161_));
  NAND2_X1  g0719(.A1(new_n1096_), .A2(new_n1098_), .ZN(new_n1162_));
  NAND2_X1  g0720(.A1(new_n1111_), .A2(new_n1113_), .ZN(new_n1163_));
  OAI211_X1 g0721(.A(new_n1161_), .B(new_n1162_), .C1(new_n1109_), .C2(new_n1163_), .ZN(new_n1164_));
  OAI21_X1  g0722(.A(new_n1104_), .B1(new_n1160_), .B2(new_n1164_), .ZN(new_n1165_));
  INV_X1    g0723(.A(new_n1048_), .ZN(new_n1166_));
  OR3_X1    g0724(.A1(new_n1165_), .A2(new_n1092_), .A3(new_n1166_), .ZN(new_n1167_));
  NOR2_X1   g0725(.A1(new_n1009_), .A2(new_n662_), .ZN(new_n1168_));
  XNOR2_X1  g0726(.A(new_n1002_), .B(KEYINPUT49), .ZN(new_n1169_));
  NAND2_X1  g0727(.A1(new_n1169_), .A2(new_n509_), .ZN(new_n1170_));
  INV_X1    g0728(.A(new_n992_), .ZN(new_n1171_));
  OAI22_X1  g0729(.A1(new_n1000_), .A2(new_n1170_), .B1(new_n1171_), .B2(new_n996_), .ZN(new_n1172_));
  NAND4_X1  g0730(.A1(new_n984_), .A2(new_n986_), .A3(new_n987_), .A4(new_n1172_), .ZN(new_n1173_));
  INV_X1    g0731(.A(new_n1173_), .ZN(new_n1174_));
  OR2_X1    g0732(.A1(new_n1174_), .A2(KEYINPUT50), .ZN(new_n1175_));
  NAND2_X1  g0733(.A1(new_n1174_), .A2(KEYINPUT50), .ZN(new_n1176_));
  INV_X1    g0734(.A(new_n991_), .ZN(new_n1177_));
  NAND3_X1  g0735(.A1(new_n987_), .A2(new_n1177_), .A3(new_n990_), .ZN(new_n1178_));
  AND2_X1   g0736(.A1(new_n984_), .A2(new_n1178_), .ZN(new_n1179_));
  OAI211_X1 g0737(.A(new_n1175_), .B(new_n1176_), .C1(new_n985_), .C2(new_n1179_), .ZN(new_n1180_));
  AOI21_X1  g0738(.A(new_n1168_), .B1(new_n1180_), .B2(new_n1013_), .ZN(new_n1181_));
  NAND4_X1  g0739(.A1(new_n1016_), .A2(new_n1094_), .A3(new_n1167_), .A4(new_n1181_), .ZN(G258));
  NAND4_X1  g0740(.A1(new_n1016_), .A2(new_n1094_), .A3(new_n1167_), .A4(new_n1181_), .ZN(G264));
  AOI21_X1  g0741(.A(new_n686_), .B1(new_n615_), .B2(new_n667_), .ZN(new_n1184_));
  INV_X1    g0742(.A(new_n823_), .ZN(new_n1185_));
  NOR2_X1   g0743(.A1(new_n842_), .A2(new_n1185_), .ZN(new_n1186_));
  NOR2_X1   g0744(.A1(new_n768_), .A2(new_n748_), .ZN(new_n1187_));
  INV_X1    g0745(.A(new_n802_), .ZN(new_n1188_));
  NAND2_X1  g0746(.A1(new_n808_), .A2(KEYINPUT54), .ZN(new_n1189_));
  OR3_X1    g0747(.A1(new_n805_), .A2(KEYINPUT54), .A3(G4405), .ZN(new_n1190_));
  AND3_X1   g0748(.A1(new_n1189_), .A2(new_n1190_), .A3(new_n809_), .ZN(new_n1191_));
  INV_X1    g0749(.A(new_n814_), .ZN(new_n1192_));
  NOR3_X1   g0750(.A1(new_n1188_), .A2(new_n1191_), .A3(new_n1192_), .ZN(new_n1193_));
  INV_X1    g0751(.A(new_n862_), .ZN(new_n1194_));
  NAND4_X1  g0752(.A1(new_n1187_), .A2(new_n1193_), .A3(G4526), .A4(new_n1194_), .ZN(new_n1195_));
  AND2_X1   g0753(.A1(new_n739_), .A2(KEYINPUT55), .ZN(new_n1196_));
  NOR2_X1   g0754(.A1(new_n739_), .A2(KEYINPUT55), .ZN(new_n1197_));
  NOR3_X1   g0755(.A1(new_n1195_), .A2(new_n1196_), .A3(new_n1197_), .ZN(new_n1198_));
  OAI21_X1  g0756(.A(new_n1186_), .B1(new_n1198_), .B2(new_n865_), .ZN(new_n1199_));
  NAND3_X1  g0757(.A1(new_n1199_), .A2(new_n840_), .A3(new_n875_), .ZN(new_n1200_));
  AND2_X1   g0758(.A1(new_n1193_), .A2(new_n1194_), .ZN(new_n1201_));
  NAND2_X1  g0759(.A1(new_n1201_), .A2(new_n1186_), .ZN(new_n1202_));
  INV_X1    g0760(.A(new_n1187_), .ZN(new_n1203_));
  OAI21_X1  g0761(.A(new_n777_), .B1(new_n734_), .B2(new_n1203_), .ZN(new_n1204_));
  INV_X1    g0762(.A(KEYINPUT53), .ZN(new_n1205_));
  AOI21_X1  g0763(.A(new_n1202_), .B1(new_n1204_), .B2(new_n1205_), .ZN(new_n1206_));
  OAI211_X1 g0764(.A(new_n777_), .B(KEYINPUT53), .C1(new_n734_), .C2(new_n1203_), .ZN(new_n1207_));
  AOI21_X1  g0765(.A(new_n1200_), .B1(new_n1206_), .B2(new_n1207_), .ZN(new_n1208_));
  OAI21_X1  g0766(.A(new_n1184_), .B1(new_n1208_), .B2(new_n895_), .ZN(G270));
  INV_X1    g0767(.A(new_n504_), .ZN(new_n1210_));
  NAND2_X1  g0768(.A1(new_n716_), .A2(new_n718_), .ZN(new_n1211_));
  NOR3_X1   g0769(.A1(new_n735_), .A2(new_n505_), .A3(new_n1211_), .ZN(new_n1212_));
  AOI21_X1  g0770(.A(new_n1210_), .B1(new_n1212_), .B2(KEYINPUT56), .ZN(new_n1213_));
  OAI21_X1  g0771(.A(new_n1213_), .B1(KEYINPUT56), .B2(new_n1212_), .ZN(new_n1214_));
  INV_X1    g0772(.A(new_n732_), .ZN(new_n1215_));
  NAND2_X1  g0773(.A1(new_n1214_), .A2(new_n1215_), .ZN(new_n1216_));
  INV_X1    g0774(.A(new_n737_), .ZN(new_n1217_));
  XNOR2_X1  g0775(.A(new_n1216_), .B(new_n1217_), .ZN(new_n1218_));
  XNOR2_X1  g0776(.A(KEYINPUT57), .B(KEYINPUT58), .ZN(new_n1219_));
  XNOR2_X1  g0777(.A(new_n1218_), .B(new_n1219_), .ZN(G388));
  XNOR2_X1  g0778(.A(new_n702_), .B(KEYINPUT59), .ZN(new_n1221_));
  OAI21_X1  g0779(.A(new_n1221_), .B1(new_n723_), .B2(new_n705_), .ZN(new_n1222_));
  INV_X1    g0780(.A(new_n1211_), .ZN(new_n1223_));
  NAND2_X1  g0781(.A1(new_n709_), .A2(new_n1223_), .ZN(new_n1224_));
  INV_X1    g0782(.A(new_n1224_), .ZN(new_n1225_));
  INV_X1    g0783(.A(new_n501_), .ZN(new_n1226_));
  OAI21_X1  g0784(.A(new_n1226_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n1227_));
  AOI21_X1  g0785(.A(new_n1222_), .B1(new_n1225_), .B2(new_n1227_), .ZN(new_n1228_));
  XNOR2_X1  g0786(.A(new_n1228_), .B(KEYINPUT60), .ZN(new_n1229_));
  XNOR2_X1  g0787(.A(new_n1229_), .B(new_n731_), .ZN(G391));
  AOI21_X1  g0788(.A(new_n715_), .B1(new_n714_), .B2(KEYINPUT62), .ZN(new_n1231_));
  OAI21_X1  g0789(.A(new_n1231_), .B1(KEYINPUT62), .B2(new_n714_), .ZN(new_n1232_));
  XOR2_X1   g0790(.A(KEYINPUT14), .B(G3705), .Z(new_n1233_));
  AOI21_X1  g0791(.A(new_n1233_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n1234_));
  AOI21_X1  g0792(.A(new_n1226_), .B1(new_n1234_), .B2(KEYINPUT62), .ZN(new_n1235_));
  AND2_X1   g0793(.A1(new_n1232_), .A2(new_n1235_), .ZN(new_n1236_));
  INV_X1    g0794(.A(new_n1236_), .ZN(new_n1237_));
  INV_X1    g0795(.A(new_n738_), .ZN(new_n1238_));
  INV_X1    g0796(.A(KEYINPUT61), .ZN(new_n1239_));
  AOI22_X1  g0797(.A1(new_n1238_), .A2(G4526), .B1(new_n1239_), .B2(new_n723_), .ZN(new_n1240_));
  OAI211_X1 g0798(.A(new_n1237_), .B(new_n1240_), .C1(new_n1239_), .C2(new_n723_), .ZN(new_n1241_));
  XNOR2_X1  g0799(.A(new_n705_), .B(KEYINPUT63), .ZN(new_n1242_));
  XNOR2_X1  g0800(.A(new_n1241_), .B(new_n1242_), .ZN(G394));
  XNOR2_X1  g0801(.A(new_n1211_), .B(new_n1227_), .ZN(G397));
  INV_X1    g0802(.A(new_n760_), .ZN(new_n1245_));
  OAI21_X1  g0803(.A(new_n759_), .B1(new_n753_), .B2(new_n1245_), .ZN(new_n1246_));
  INV_X1    g0804(.A(new_n1246_), .ZN(new_n1247_));
  OAI21_X1  g0805(.A(new_n774_), .B1(new_n1247_), .B2(new_n748_), .ZN(new_n1248_));
  NAND2_X1  g0806(.A1(new_n741_), .A2(new_n1248_), .ZN(new_n1249_));
  XOR2_X1   g0807(.A(new_n772_), .B(KEYINPUT64), .Z(new_n1250_));
  NOR2_X1   g0808(.A1(new_n1250_), .A2(new_n775_), .ZN(new_n1251_));
  XOR2_X1   g0809(.A(new_n1251_), .B(KEYINPUT65), .Z(new_n1252_));
  OAI21_X1  g0810(.A(new_n1249_), .B1(new_n1252_), .B2(new_n741_), .ZN(new_n1253_));
  NAND2_X1  g0811(.A1(new_n766_), .A2(new_n767_), .ZN(new_n1254_));
  XNOR2_X1  g0812(.A(new_n1253_), .B(new_n1254_), .ZN(G376));
  INV_X1    g0813(.A(new_n771_), .ZN(new_n1256_));
  NOR2_X1   g0814(.A1(new_n1256_), .A2(new_n770_), .ZN(new_n1257_));
  XOR2_X1   g0815(.A(new_n749_), .B(new_n1257_), .Z(new_n1258_));
  NAND2_X1  g0816(.A1(new_n742_), .A2(new_n1258_), .ZN(new_n1259_));
  INV_X1    g0817(.A(new_n748_), .ZN(new_n1260_));
  XNOR2_X1  g0818(.A(new_n1246_), .B(new_n1260_), .ZN(new_n1261_));
  OAI21_X1  g0819(.A(new_n1259_), .B1(new_n742_), .B2(new_n1261_), .ZN(G379));
  AOI21_X1  g0820(.A(new_n754_), .B1(new_n741_), .B2(new_n752_), .ZN(new_n1263_));
  XNOR2_X1  g0821(.A(new_n1263_), .B(new_n762_), .ZN(G382));
  XOR2_X1   g0822(.A(new_n755_), .B(KEYINPUT66), .Z(new_n1265_));
  XNOR2_X1  g0823(.A(new_n741_), .B(new_n1265_), .ZN(G385));
  XOR2_X1   g0824(.A(new_n805_), .B(new_n797_), .Z(new_n1267_));
  XOR2_X1   g0825(.A(new_n1267_), .B(KEYINPUT69), .Z(new_n1268_));
  XOR2_X1   g0826(.A(new_n780_), .B(new_n813_), .Z(new_n1269_));
  XNOR2_X1  g0827(.A(new_n1269_), .B(KEYINPUT68), .ZN(new_n1270_));
  NAND2_X1  g0828(.A1(new_n507_), .A2(G115), .ZN(new_n1271_));
  INV_X1    g0829(.A(G227), .ZN(new_n1272_));
  OAI21_X1  g0830(.A(new_n1271_), .B1(new_n507_), .B2(new_n1272_), .ZN(new_n1273_));
  XNOR2_X1  g0831(.A(new_n789_), .B(new_n1273_), .ZN(new_n1274_));
  INV_X1    g0832(.A(new_n1274_), .ZN(new_n1275_));
  NAND3_X1  g0833(.A1(new_n1268_), .A2(new_n1270_), .A3(new_n1275_), .ZN(new_n1276_));
  XNOR2_X1  g0834(.A(new_n1276_), .B(KEYINPUT70), .ZN(new_n1277_));
  OR2_X1    g0835(.A1(new_n1268_), .A2(new_n1275_), .ZN(new_n1278_));
  AOI21_X1  g0836(.A(new_n1269_), .B1(new_n1275_), .B2(new_n1267_), .ZN(new_n1279_));
  NOR2_X1   g0837(.A1(new_n1275_), .A2(new_n1267_), .ZN(new_n1280_));
  AOI22_X1  g0838(.A1(new_n1278_), .A2(new_n1279_), .B1(new_n1270_), .B2(new_n1280_), .ZN(new_n1281_));
  NAND2_X1  g0839(.A1(new_n1277_), .A2(new_n1281_), .ZN(new_n1282_));
  XOR2_X1   g0840(.A(new_n1282_), .B(new_n828_), .Z(new_n1283_));
  XNOR2_X1  g0841(.A(new_n819_), .B(KEYINPUT71), .ZN(new_n1284_));
  XNOR2_X1  g0842(.A(new_n1283_), .B(new_n1284_), .ZN(new_n1285_));
  XNOR2_X1  g0843(.A(new_n839_), .B(new_n871_), .ZN(new_n1286_));
  OR2_X1    g0844(.A1(new_n1285_), .A2(new_n1286_), .ZN(new_n1287_));
  NAND2_X1  g0845(.A1(new_n1285_), .A2(new_n1286_), .ZN(new_n1288_));
  AOI21_X1  g0846(.A(new_n536_), .B1(new_n507_), .B2(G147), .ZN(new_n1289_));
  NOR3_X1   g0847(.A1(new_n534_), .A2(KEYINPUT10), .A3(G18), .ZN(new_n1290_));
  OAI21_X1  g0848(.A(new_n539_), .B1(new_n1289_), .B2(new_n1290_), .ZN(new_n1291_));
  NAND2_X1  g0849(.A1(new_n507_), .A2(G141), .ZN(new_n1292_));
  INV_X1    g0850(.A(G161), .ZN(new_n1293_));
  OAI21_X1  g0851(.A(new_n1292_), .B1(new_n507_), .B2(new_n1293_), .ZN(new_n1294_));
  XNOR2_X1  g0852(.A(new_n1291_), .B(new_n1294_), .ZN(new_n1295_));
  XNOR2_X1  g0853(.A(new_n1295_), .B(new_n524_), .ZN(new_n1296_));
  NAND2_X1  g0854(.A1(new_n575_), .A2(new_n508_), .ZN(new_n1297_));
  OAI21_X1  g0855(.A(new_n1297_), .B1(new_n511_), .B2(new_n575_), .ZN(new_n1298_));
  XNOR2_X1  g0856(.A(new_n1296_), .B(new_n1298_), .ZN(new_n1299_));
  XOR2_X1   g0857(.A(new_n567_), .B(new_n517_), .Z(new_n1300_));
  XNOR2_X1  g0858(.A(new_n1299_), .B(new_n1300_), .ZN(new_n1301_));
  OR3_X1    g0859(.A1(new_n592_), .A2(new_n507_), .A3(G155), .ZN(new_n1302_));
  OAI21_X1  g0860(.A(new_n1302_), .B1(new_n582_), .B2(new_n591_), .ZN(new_n1303_));
  XOR2_X1   g0861(.A(new_n1303_), .B(new_n602_), .Z(new_n1304_));
  AND2_X1   g0862(.A1(new_n1301_), .A2(new_n1304_), .ZN(new_n1305_));
  NOR2_X1   g0863(.A1(new_n1301_), .A2(new_n1304_), .ZN(new_n1306_));
  OAI21_X1  g0864(.A(new_n641_), .B1(new_n507_), .B2(G215), .ZN(new_n1307_));
  OAI21_X1  g0865(.A(new_n1307_), .B1(new_n625_), .B2(new_n641_), .ZN(new_n1308_));
  OAI22_X1  g0866(.A1(new_n648_), .A2(new_n617_), .B1(new_n649_), .B2(new_n616_), .ZN(new_n1309_));
  XNOR2_X1  g0867(.A(new_n1308_), .B(new_n1309_), .ZN(new_n1310_));
  NOR2_X1   g0868(.A1(new_n1310_), .A2(KEYINPUT67), .ZN(new_n1311_));
  XNOR2_X1  g0869(.A(G211), .B(G212), .ZN(new_n1312_));
  XNOR2_X1  g0870(.A(new_n1312_), .B(new_n633_), .ZN(new_n1313_));
  NAND3_X1  g0871(.A1(new_n1313_), .A2(G18), .A3(new_n509_), .ZN(new_n1314_));
  XNOR2_X1  g0872(.A(new_n1311_), .B(new_n1314_), .ZN(new_n1315_));
  NAND2_X1  g0873(.A1(new_n507_), .A2(G41), .ZN(new_n1316_));
  INV_X1    g0874(.A(G229), .ZN(new_n1317_));
  OAI21_X1  g0875(.A(new_n1316_), .B1(new_n507_), .B2(new_n1317_), .ZN(new_n1318_));
  XNOR2_X1  g0876(.A(new_n751_), .B(new_n1318_), .ZN(new_n1319_));
  XNOR2_X1  g0877(.A(new_n1319_), .B(new_n695_), .ZN(new_n1320_));
  NAND2_X1  g0878(.A1(new_n507_), .A2(G44), .ZN(new_n1321_));
  INV_X1    g0879(.A(G239), .ZN(new_n1322_));
  OAI21_X1  g0880(.A(new_n1321_), .B1(new_n507_), .B2(new_n1322_), .ZN(new_n1323_));
  XNOR2_X1  g0881(.A(new_n1323_), .B(new_n700_), .ZN(new_n1324_));
  XNOR2_X1  g0882(.A(new_n1324_), .B(new_n691_), .ZN(new_n1325_));
  XOR2_X1   g0883(.A(new_n1320_), .B(new_n1325_), .Z(new_n1326_));
  XNOR2_X1  g0884(.A(new_n714_), .B(new_n745_), .ZN(new_n1327_));
  XNOR2_X1  g0885(.A(new_n765_), .B(new_n758_), .ZN(new_n1328_));
  XNOR2_X1  g0886(.A(new_n1327_), .B(new_n1328_), .ZN(new_n1329_));
  INV_X1    g0887(.A(new_n1329_), .ZN(new_n1330_));
  OAI21_X1  g0888(.A(new_n1315_), .B1(new_n1326_), .B2(new_n1330_), .ZN(new_n1331_));
  INV_X1    g0889(.A(new_n1326_), .ZN(new_n1332_));
  NOR2_X1   g0890(.A1(new_n1332_), .A2(new_n1329_), .ZN(new_n1333_));
  NOR4_X1   g0891(.A1(new_n1305_), .A2(new_n1306_), .A3(new_n1331_), .A4(new_n1333_), .ZN(new_n1334_));
  NAND3_X1  g0892(.A1(new_n1287_), .A2(new_n1288_), .A3(new_n1334_), .ZN(G412));
  XNOR2_X1  g0893(.A(new_n975_), .B(new_n983_), .ZN(new_n1336_));
  XOR2_X1   g0894(.A(new_n990_), .B(new_n994_), .Z(new_n1337_));
  NAND2_X1  g0895(.A1(new_n1336_), .A2(new_n1337_), .ZN(new_n1338_));
  NAND2_X1  g0896(.A1(new_n507_), .A2(G114), .ZN(new_n1339_));
  OAI21_X1  g0897(.A(new_n1339_), .B1(new_n507_), .B2(G1459), .ZN(new_n1340_));
  XNOR2_X1  g0898(.A(new_n1169_), .B(new_n1340_), .ZN(new_n1341_));
  NOR2_X1   g0899(.A1(new_n1338_), .A2(new_n1341_), .ZN(new_n1342_));
  XOR2_X1   g0900(.A(new_n1342_), .B(KEYINPUT73), .Z(new_n1343_));
  OR2_X1    g0901(.A1(new_n1336_), .A2(new_n1337_), .ZN(new_n1344_));
  NAND3_X1  g0902(.A1(new_n1344_), .A2(new_n1338_), .A3(new_n1341_), .ZN(new_n1345_));
  OAI21_X1  g0903(.A(new_n1345_), .B1(new_n1341_), .B2(new_n1344_), .ZN(new_n1346_));
  NOR2_X1   g0904(.A1(new_n1343_), .A2(new_n1346_), .ZN(new_n1347_));
  MUX2_X1   g0905(.A(new_n1005_), .B(G1492), .S(G18), .Z(new_n1348_));
  XNOR2_X1  g0906(.A(new_n1347_), .B(new_n1348_), .ZN(new_n1349_));
  MUX2_X1   g0907(.A(new_n1010_), .B(G1496), .S(G18), .Z(new_n1350_));
  XNOR2_X1  g0908(.A(new_n1349_), .B(new_n1350_), .ZN(new_n1351_));
  NOR2_X1   g0909(.A1(new_n507_), .A2(G3698), .ZN(new_n1352_));
  AOI21_X1  g0910(.A(new_n1352_), .B1(new_n507_), .B2(G69), .ZN(new_n1353_));
  XNOR2_X1  g0911(.A(new_n1353_), .B(new_n1141_), .ZN(new_n1354_));
  XNOR2_X1  g0912(.A(new_n1354_), .B(new_n1108_), .ZN(new_n1355_));
  XNOR2_X1  g0913(.A(new_n1355_), .B(new_n1113_), .ZN(new_n1356_));
  XNOR2_X1  g0914(.A(new_n1356_), .B(new_n1098_), .ZN(new_n1357_));
  XNOR2_X1  g0915(.A(new_n1357_), .B(new_n1125_), .ZN(new_n1358_));
  NAND2_X1  g0916(.A1(G18), .A2(G3701), .ZN(new_n1359_));
  OAI21_X1  g0917(.A(new_n1359_), .B1(G18), .B2(G70), .ZN(new_n1360_));
  XNOR2_X1  g0918(.A(new_n1132_), .B(new_n1360_), .ZN(new_n1361_));
  XNOR2_X1  g0919(.A(new_n1361_), .B(new_n1137_), .ZN(new_n1362_));
  XNOR2_X1  g0920(.A(new_n1362_), .B(new_n1119_), .ZN(new_n1363_));
  XNOR2_X1  g0921(.A(new_n1358_), .B(new_n1363_), .ZN(new_n1364_));
  NOR2_X1   g0922(.A1(new_n1351_), .A2(new_n1364_), .ZN(new_n1365_));
  XNOR2_X1  g0923(.A(new_n960_), .B(new_n950_), .ZN(new_n1366_));
  XNOR2_X1  g0924(.A(new_n1366_), .B(new_n941_), .ZN(new_n1367_));
  NOR2_X1   g0925(.A1(G18), .A2(G82), .ZN(new_n1368_));
  AOI21_X1  g0926(.A(new_n1368_), .B1(G18), .B2(G2208), .ZN(new_n1369_));
  INV_X1    g0927(.A(new_n1369_), .ZN(new_n1370_));
  NAND2_X1  g0928(.A1(new_n1367_), .A2(new_n1370_), .ZN(new_n1371_));
  XNOR2_X1  g0929(.A(new_n1366_), .B(new_n940_), .ZN(new_n1372_));
  NAND2_X1  g0930(.A1(new_n1372_), .A2(new_n1369_), .ZN(new_n1373_));
  NAND3_X1  g0931(.A1(new_n1371_), .A2(new_n1373_), .A3(KEYINPUT72), .ZN(new_n1374_));
  XNOR2_X1  g0932(.A(new_n1374_), .B(new_n922_), .ZN(new_n1375_));
  XNOR2_X1  g0933(.A(new_n1375_), .B(new_n907_), .ZN(new_n1376_));
  XNOR2_X1  g0934(.A(new_n901_), .B(new_n926_), .ZN(new_n1377_));
  XNOR2_X1  g0935(.A(new_n1377_), .B(new_n932_), .ZN(new_n1378_));
  XNOR2_X1  g0936(.A(new_n1378_), .B(new_n915_), .ZN(new_n1379_));
  XNOR2_X1  g0937(.A(new_n1376_), .B(new_n1379_), .ZN(new_n1380_));
  XNOR2_X1  g0938(.A(new_n1070_), .B(new_n1076_), .ZN(new_n1381_));
  XNOR2_X1  g0939(.A(new_n1381_), .B(new_n1066_), .ZN(new_n1382_));
  XNOR2_X1  g0940(.A(new_n1382_), .B(new_n1061_), .ZN(new_n1383_));
  XNOR2_X1  g0941(.A(new_n1032_), .B(new_n1026_), .ZN(new_n1384_));
  XNOR2_X1  g0942(.A(new_n1383_), .B(new_n1384_), .ZN(new_n1385_));
  NOR2_X1   g0943(.A1(G18), .A2(G58), .ZN(new_n1386_));
  AOI21_X1  g0944(.A(new_n1386_), .B1(G18), .B2(G4393), .ZN(new_n1387_));
  XNOR2_X1  g0945(.A(new_n1038_), .B(new_n1387_), .ZN(new_n1388_));
  XNOR2_X1  g0946(.A(new_n1385_), .B(new_n1388_), .ZN(new_n1389_));
  XOR2_X1   g0947(.A(new_n1020_), .B(new_n1050_), .Z(new_n1390_));
  XNOR2_X1  g0948(.A(new_n1389_), .B(new_n1390_), .ZN(new_n1391_));
  NAND3_X1  g0949(.A1(new_n1365_), .A2(new_n1380_), .A3(new_n1391_), .ZN(new_n1392_));
  NAND2_X1  g0950(.A1(new_n1392_), .A2(KEYINPUT74), .ZN(new_n1393_));
  INV_X1    g0951(.A(KEYINPUT74), .ZN(new_n1394_));
  NAND4_X1  g0952(.A1(new_n1365_), .A2(new_n1380_), .A3(new_n1394_), .A4(new_n1391_), .ZN(new_n1395_));
  NAND2_X1  g0953(.A1(new_n1393_), .A2(new_n1395_), .ZN(G414));
  INV_X1    g0954(.A(G198), .ZN(new_n1397_));
  OAI21_X1  g0955(.A(new_n1316_), .B1(new_n507_), .B2(new_n1397_), .ZN(new_n1398_));
  INV_X1    g0956(.A(G208), .ZN(new_n1399_));
  OAI21_X1  g0957(.A(new_n1321_), .B1(new_n507_), .B2(new_n1399_), .ZN(new_n1400_));
  XOR2_X1   g0958(.A(new_n1398_), .B(new_n1400_), .Z(new_n1401_));
  XNOR2_X1  g0959(.A(new_n1129_), .B(new_n1117_), .ZN(new_n1402_));
  OR2_X1    g0960(.A1(new_n1401_), .A2(new_n1402_), .ZN(new_n1403_));
  XOR2_X1   g0961(.A(new_n1135_), .B(new_n1139_), .Z(new_n1404_));
  NOR2_X1   g0962(.A1(new_n1403_), .A2(new_n1404_), .ZN(new_n1405_));
  XOR2_X1   g0963(.A(new_n1405_), .B(KEYINPUT76), .Z(new_n1406_));
  NAND2_X1  g0964(.A1(new_n1401_), .A2(new_n1402_), .ZN(new_n1407_));
  NOR2_X1   g0965(.A1(new_n1407_), .A2(new_n1404_), .ZN(new_n1408_));
  XOR2_X1   g0966(.A(new_n1408_), .B(KEYINPUT75), .Z(new_n1409_));
  NAND3_X1  g0967(.A1(new_n1403_), .A2(new_n1404_), .A3(new_n1407_), .ZN(new_n1410_));
  NAND3_X1  g0968(.A1(new_n1406_), .A2(new_n1409_), .A3(new_n1410_), .ZN(new_n1411_));
  XOR2_X1   g0969(.A(new_n1096_), .B(KEYINPUT77), .Z(new_n1412_));
  XNOR2_X1  g0970(.A(new_n1411_), .B(new_n1412_), .ZN(new_n1413_));
  XOR2_X1   g0971(.A(new_n1111_), .B(new_n1106_), .Z(new_n1414_));
  XNOR2_X1  g0972(.A(new_n1414_), .B(new_n1122_), .ZN(new_n1415_));
  XNOR2_X1  g0973(.A(new_n1413_), .B(new_n1415_), .ZN(new_n1416_));
  NAND2_X1  g0974(.A1(new_n920_), .A2(new_n911_), .ZN(new_n1417_));
  OAI21_X1  g0975(.A(new_n1417_), .B1(new_n913_), .B2(new_n920_), .ZN(new_n1418_));
  XNOR2_X1  g0976(.A(new_n1418_), .B(new_n898_), .ZN(new_n1419_));
  XNOR2_X1  g0977(.A(new_n1419_), .B(new_n927_), .ZN(new_n1420_));
  INV_X1    g0978(.A(G181), .ZN(new_n1421_));
  OAI21_X1  g0979(.A(new_n1292_), .B1(new_n507_), .B2(new_n1421_), .ZN(new_n1422_));
  XNOR2_X1  g0980(.A(new_n1422_), .B(new_n904_), .ZN(new_n1423_));
  XNOR2_X1  g0981(.A(new_n1423_), .B(new_n947_), .ZN(new_n1424_));
  XNOR2_X1  g0982(.A(new_n1424_), .B(new_n962_), .ZN(new_n1425_));
  XNOR2_X1  g0983(.A(new_n1420_), .B(new_n1425_), .ZN(new_n1426_));
  XOR2_X1   g0984(.A(new_n936_), .B(new_n930_), .Z(new_n1427_));
  XNOR2_X1  g0985(.A(new_n1426_), .B(new_n1427_), .ZN(new_n1428_));
  INV_X1    g0986(.A(G197), .ZN(new_n1429_));
  OAI21_X1  g0987(.A(new_n1271_), .B1(new_n507_), .B2(new_n1429_), .ZN(new_n1430_));
  XOR2_X1   g0988(.A(new_n1074_), .B(new_n1430_), .Z(new_n1431_));
  XNOR2_X1  g0989(.A(new_n1431_), .B(new_n1064_), .ZN(new_n1432_));
  XOR2_X1   g0990(.A(new_n1024_), .B(new_n1053_), .Z(new_n1433_));
  XNOR2_X1  g0991(.A(new_n1432_), .B(new_n1433_), .ZN(new_n1434_));
  XOR2_X1   g0992(.A(new_n1072_), .B(KEYINPUT78), .Z(new_n1435_));
  XOR2_X1   g0993(.A(new_n1435_), .B(new_n1057_), .Z(new_n1436_));
  XNOR2_X1  g0994(.A(new_n1434_), .B(new_n1436_), .ZN(new_n1437_));
  XNOR2_X1  g0995(.A(new_n1030_), .B(new_n1039_), .ZN(new_n1438_));
  XNOR2_X1  g0996(.A(new_n1018_), .B(KEYINPUT79), .ZN(new_n1439_));
  XNOR2_X1  g0997(.A(new_n1438_), .B(new_n1439_), .ZN(new_n1440_));
  AND2_X1   g0998(.A1(new_n1437_), .A2(new_n1440_), .ZN(new_n1441_));
  NOR2_X1   g0999(.A1(new_n1437_), .A2(new_n1440_), .ZN(new_n1442_));
  MUX2_X1   g1000(.A(new_n976_), .B(new_n977_), .S(new_n979_), .Z(new_n1443_));
  MUX2_X1   g1001(.A(new_n995_), .B(new_n998_), .S(new_n991_), .Z(new_n1444_));
  XNOR2_X1  g1002(.A(new_n1443_), .B(new_n1444_), .ZN(new_n1445_));
  NOR3_X1   g1003(.A1(new_n573_), .A2(new_n507_), .A3(G170), .ZN(new_n1446_));
  XNOR2_X1  g1004(.A(new_n1446_), .B(KEYINPUT80), .ZN(new_n1447_));
  XNOR2_X1  g1005(.A(new_n1445_), .B(new_n1447_), .ZN(new_n1448_));
  INV_X1    g1006(.A(G164), .ZN(new_n1449_));
  OR2_X1    g1007(.A1(new_n1449_), .A2(G165), .ZN(new_n1450_));
  NAND2_X1  g1008(.A1(new_n1449_), .A2(G165), .ZN(new_n1451_));
  AOI211_X1 g1009(.A(new_n507_), .B(new_n573_), .C1(new_n1450_), .C2(new_n1451_), .ZN(new_n1452_));
  XNOR2_X1  g1010(.A(new_n1448_), .B(new_n1452_), .ZN(new_n1453_));
  NOR3_X1   g1011(.A1(new_n1441_), .A2(new_n1442_), .A3(new_n1453_), .ZN(new_n1454_));
  NAND3_X1  g1012(.A1(new_n1416_), .A2(new_n1428_), .A3(new_n1454_), .ZN(G416));
  NAND2_X1  g1013(.A1(new_n1165_), .A2(new_n1086_), .ZN(new_n1456_));
  AOI21_X1  g1014(.A(new_n1043_), .B1(new_n1456_), .B2(new_n1048_), .ZN(new_n1457_));
  OAI21_X1  g1015(.A(new_n972_), .B1(new_n1457_), .B2(new_n1091_), .ZN(new_n1458_));
  AOI21_X1  g1016(.A(new_n1180_), .B1(new_n1458_), .B2(new_n1004_), .ZN(new_n1459_));
  OAI22_X1  g1017(.A1(new_n1459_), .A2(new_n1012_), .B1(new_n662_), .B2(new_n1009_), .ZN(new_n1460_));
  XNOR2_X1  g1018(.A(new_n1460_), .B(KEYINPUT81), .ZN(G249));
  NOR2_X1   g1019(.A1(new_n888_), .A2(new_n540_), .ZN(new_n1462_));
  XNOR2_X1  g1020(.A(new_n878_), .B(new_n1462_), .ZN(G295));
  NOR2_X1   g1021(.A1(new_n878_), .A2(new_n893_), .ZN(new_n1464_));
  NOR2_X1   g1022(.A1(new_n1464_), .A2(new_n615_), .ZN(new_n1465_));
  NAND2_X1  g1023(.A1(new_n1465_), .A2(new_n639_), .ZN(new_n1466_));
  INV_X1    g1024(.A(new_n639_), .ZN(new_n1467_));
  OAI21_X1  g1025(.A(new_n1467_), .B1(new_n1464_), .B2(new_n615_), .ZN(new_n1468_));
  NAND2_X1  g1026(.A1(new_n1466_), .A2(new_n1468_), .ZN(new_n1469_));
  XOR2_X1   g1027(.A(new_n1469_), .B(KEYINPUT82), .Z(G324));
  XNOR2_X1  g1028(.A(new_n1457_), .B(KEYINPUT83), .ZN(G252));
  AND3_X1   g1029(.A1(new_n1204_), .A2(new_n1186_), .A3(new_n1201_), .ZN(new_n1472_));
  OAI21_X1  g1030(.A(new_n894_), .B1(new_n1472_), .B2(new_n1200_), .ZN(new_n1473_));
  XNOR2_X1  g1031(.A(new_n615_), .B(KEYINPUT84), .ZN(new_n1474_));
  AND2_X1   g1032(.A1(new_n1473_), .A2(new_n1474_), .ZN(new_n1475_));
  INV_X1    g1033(.A(new_n1475_), .ZN(new_n1476_));
  AOI21_X1  g1034(.A(new_n684_), .B1(new_n1476_), .B2(new_n657_), .ZN(new_n1477_));
  OAI21_X1  g1035(.A(new_n670_), .B1(new_n1477_), .B2(new_n666_), .ZN(G276));
  INV_X1    g1036(.A(new_n527_), .ZN(new_n1479_));
  AOI21_X1  g1037(.A(KEYINPUT20), .B1(new_n517_), .B2(new_n518_), .ZN(new_n1480_));
  NOR2_X1   g1038(.A1(new_n1479_), .A2(new_n1480_), .ZN(new_n1481_));
  INV_X1    g1039(.A(new_n1481_), .ZN(new_n1482_));
  AOI21_X1  g1040(.A(new_n569_), .B1(new_n885_), .B2(new_n1482_), .ZN(new_n1483_));
  AOI21_X1  g1041(.A(new_n560_), .B1(new_n526_), .B2(new_n544_), .ZN(new_n1484_));
  INV_X1    g1042(.A(new_n1484_), .ZN(new_n1485_));
  INV_X1    g1043(.A(new_n1462_), .ZN(new_n1486_));
  NOR2_X1   g1044(.A1(new_n878_), .A2(new_n1486_), .ZN(new_n1487_));
  NAND2_X1  g1045(.A1(new_n1487_), .A2(new_n533_), .ZN(new_n1488_));
  OAI21_X1  g1046(.A(new_n543_), .B1(new_n553_), .B2(new_n559_), .ZN(new_n1489_));
  OAI211_X1 g1047(.A(new_n1483_), .B(new_n1485_), .C1(new_n1488_), .C2(new_n1489_), .ZN(new_n1490_));
  XNOR2_X1  g1048(.A(new_n1490_), .B(new_n879_), .ZN(G310));
  NOR2_X1   g1049(.A1(new_n880_), .A2(new_n889_), .ZN(new_n1492_));
  NAND2_X1  g1050(.A1(new_n1487_), .A2(new_n1492_), .ZN(new_n1493_));
  AOI21_X1  g1051(.A(new_n545_), .B1(new_n1493_), .B2(KEYINPUT85), .ZN(new_n1494_));
  OAI21_X1  g1052(.A(new_n1494_), .B1(KEYINPUT85), .B2(new_n1493_), .ZN(new_n1495_));
  XNOR2_X1  g1053(.A(new_n1495_), .B(new_n560_), .ZN(G313));
  INV_X1    g1054(.A(KEYINPUT86), .ZN(new_n1497_));
  OAI21_X1  g1055(.A(new_n1497_), .B1(new_n1479_), .B2(new_n1480_), .ZN(new_n1498_));
  NAND3_X1  g1056(.A1(new_n521_), .A2(KEYINPUT86), .A3(new_n527_), .ZN(new_n1499_));
  NAND4_X1  g1057(.A1(new_n1291_), .A2(new_n886_), .A3(new_n519_), .A4(new_n532_), .ZN(new_n1500_));
  NAND3_X1  g1058(.A1(new_n1498_), .A2(new_n1499_), .A3(new_n1500_), .ZN(new_n1501_));
  INV_X1    g1059(.A(new_n1501_), .ZN(new_n1502_));
  NAND2_X1  g1060(.A1(new_n1488_), .A2(new_n1502_), .ZN(new_n1503_));
  XNOR2_X1  g1061(.A(new_n1503_), .B(new_n880_), .ZN(G316));
  NOR2_X1   g1062(.A1(new_n1487_), .A2(new_n540_), .ZN(new_n1505_));
  XNOR2_X1  g1063(.A(new_n1505_), .B(new_n533_), .ZN(G319));
  NOR2_X1   g1064(.A1(new_n1465_), .A2(new_n647_), .ZN(new_n1507_));
  INV_X1    g1065(.A(KEYINPUT87), .ZN(new_n1508_));
  XNOR2_X1  g1066(.A(new_n638_), .B(new_n1508_), .ZN(new_n1509_));
  OAI21_X1  g1067(.A(new_n676_), .B1(new_n1509_), .B2(new_n645_), .ZN(new_n1510_));
  AOI21_X1  g1068(.A(new_n681_), .B1(new_n1510_), .B2(new_n632_), .ZN(new_n1511_));
  INV_X1    g1069(.A(new_n1511_), .ZN(new_n1512_));
  NOR2_X1   g1070(.A1(new_n1507_), .A2(new_n1512_), .ZN(new_n1513_));
  XNOR2_X1  g1071(.A(new_n1513_), .B(new_n655_), .ZN(G327));
  INV_X1    g1072(.A(new_n680_), .ZN(new_n1515_));
  NOR2_X1   g1073(.A1(new_n677_), .A2(new_n1515_), .ZN(new_n1516_));
  NAND2_X1  g1074(.A1(new_n628_), .A2(new_n630_), .ZN(new_n1517_));
  INV_X1    g1075(.A(new_n645_), .ZN(new_n1518_));
  NAND2_X1  g1076(.A1(new_n1517_), .A2(new_n1518_), .ZN(new_n1519_));
  OAI21_X1  g1077(.A(new_n1516_), .B1(new_n1468_), .B2(new_n1519_), .ZN(new_n1520_));
  XNOR2_X1  g1078(.A(new_n1520_), .B(new_n623_), .ZN(G330));
  AND2_X1   g1079(.A1(new_n1468_), .A2(new_n1509_), .ZN(new_n1522_));
  OAI211_X1 g1080(.A(new_n1517_), .B(new_n643_), .C1(new_n1522_), .C2(new_n645_), .ZN(new_n1523_));
  AOI21_X1  g1081(.A(new_n645_), .B1(new_n1468_), .B2(new_n1509_), .ZN(new_n1524_));
  INV_X1    g1082(.A(new_n643_), .ZN(new_n1525_));
  OAI21_X1  g1083(.A(new_n631_), .B1(new_n1524_), .B2(new_n1525_), .ZN(new_n1526_));
  NAND2_X1  g1084(.A1(new_n1523_), .A2(new_n1526_), .ZN(G333));
  XNOR2_X1  g1085(.A(new_n1522_), .B(new_n1518_), .ZN(G336));
  NOR4_X1   g1086(.A1(G404), .A2(G406), .A3(G408), .A4(G410), .ZN(new_n1529_));
  NOR2_X1   g1087(.A1(G412), .A2(G416), .ZN(new_n1530_));
  NAND3_X1  g1088(.A1(new_n1393_), .A2(new_n1530_), .A3(new_n1395_), .ZN(new_n1531_));
  AND2_X1   g1089(.A1(new_n1531_), .A2(KEYINPUT88), .ZN(new_n1532_));
  NOR2_X1   g1090(.A1(new_n1531_), .A2(KEYINPUT88), .ZN(new_n1533_));
  OAI21_X1  g1091(.A(new_n1529_), .B1(new_n1532_), .B2(new_n1533_), .ZN(G418));
  AOI21_X1  g1092(.A(new_n684_), .B1(new_n1507_), .B2(new_n655_), .ZN(new_n1535_));
  OAI21_X1  g1093(.A(new_n670_), .B1(new_n1535_), .B2(new_n666_), .ZN(G273));
  INV_X1    g1094(.A(new_n878_), .ZN(new_n1537_));
  AOI21_X1  g1095(.A(new_n572_), .B1(new_n1537_), .B2(new_n892_), .ZN(new_n1538_));
  INV_X1    g1096(.A(new_n1538_), .ZN(new_n1539_));
  OAI21_X1  g1097(.A(new_n578_), .B1(new_n595_), .B2(new_n610_), .ZN(new_n1540_));
  NAND2_X1  g1098(.A1(new_n1539_), .A2(new_n1540_), .ZN(new_n1541_));
  NAND2_X1  g1099(.A1(new_n611_), .A2(new_n612_), .ZN(new_n1542_));
  NAND2_X1  g1100(.A1(new_n1542_), .A2(new_n578_), .ZN(new_n1543_));
  NAND2_X1  g1101(.A1(new_n1538_), .A2(new_n1543_), .ZN(new_n1544_));
  NAND2_X1  g1102(.A1(new_n1541_), .A2(new_n1544_), .ZN(new_n1545_));
  INV_X1    g1103(.A(new_n605_), .ZN(new_n1546_));
  XNOR2_X1  g1104(.A(new_n1545_), .B(new_n1546_), .ZN(G298));
  NAND2_X1  g1105(.A1(new_n612_), .A2(new_n609_), .ZN(new_n1548_));
  XNOR2_X1  g1106(.A(new_n581_), .B(new_n1548_), .ZN(new_n1549_));
  NAND2_X1  g1107(.A1(new_n1538_), .A2(new_n1549_), .ZN(new_n1550_));
  XOR2_X1   g1108(.A(new_n580_), .B(KEYINPUT89), .Z(new_n1551_));
  NAND2_X1  g1109(.A1(new_n596_), .A2(new_n609_), .ZN(new_n1552_));
  XOR2_X1   g1110(.A(new_n1551_), .B(new_n1552_), .Z(new_n1553_));
  OAI21_X1  g1111(.A(new_n1550_), .B1(new_n1538_), .B2(new_n1553_), .ZN(new_n1554_));
  XOR2_X1   g1112(.A(new_n1554_), .B(KEYINPUT90), .Z(G301));
  XNOR2_X1  g1113(.A(new_n589_), .B(new_n600_), .ZN(new_n1556_));
  XNOR2_X1  g1114(.A(new_n1556_), .B(KEYINPUT91), .ZN(new_n1557_));
  NAND2_X1  g1115(.A1(new_n1538_), .A2(new_n1557_), .ZN(new_n1558_));
  XNOR2_X1  g1116(.A(new_n589_), .B(new_n594_), .ZN(new_n1559_));
  OAI21_X1  g1117(.A(new_n1558_), .B1(new_n1538_), .B2(new_n1559_), .ZN(G304));
  NAND2_X1  g1118(.A1(new_n599_), .A2(new_n593_), .ZN(new_n1561_));
  XOR2_X1   g1119(.A(new_n1538_), .B(new_n1561_), .Z(G307));
  INV_X1    g1120(.A(new_n794_), .ZN(new_n1563_));
  XNOR2_X1  g1121(.A(new_n779_), .B(new_n1563_), .ZN(G344));
  NAND2_X1  g1122(.A1(new_n1507_), .A2(new_n655_), .ZN(new_n1565_));
  NAND2_X1  g1123(.A1(new_n1565_), .A2(new_n685_), .ZN(new_n1566_));
  AND2_X1   g1124(.A1(new_n661_), .A2(new_n663_), .ZN(new_n1567_));
  NAND2_X1  g1125(.A1(new_n664_), .A2(G38), .ZN(new_n1568_));
  AOI22_X1  g1126(.A1(new_n1567_), .A2(new_n1568_), .B1(G1496), .B2(new_n660_), .ZN(new_n1569_));
  NAND2_X1  g1127(.A1(new_n1566_), .A2(new_n1569_), .ZN(new_n1570_));
  INV_X1    g1128(.A(new_n1568_), .ZN(new_n1571_));
  AOI22_X1  g1129(.A1(new_n659_), .A2(new_n1571_), .B1(new_n665_), .B2(new_n663_), .ZN(new_n1572_));
  XNOR2_X1  g1130(.A(new_n1572_), .B(KEYINPUT92), .ZN(new_n1573_));
  NAND2_X1  g1131(.A1(new_n1535_), .A2(new_n1573_), .ZN(new_n1574_));
  NAND2_X1  g1132(.A1(new_n1570_), .A2(new_n1574_), .ZN(G422));
  NAND2_X1  g1133(.A1(new_n1570_), .A2(new_n1574_), .ZN(G469));
  NAND2_X1  g1134(.A1(new_n659_), .A2(G38), .ZN(new_n1577_));
  NAND2_X1  g1135(.A1(new_n661_), .A2(new_n1577_), .ZN(new_n1578_));
  NAND2_X1  g1136(.A1(new_n1566_), .A2(new_n1578_), .ZN(new_n1579_));
  NAND3_X1  g1137(.A1(new_n1535_), .A2(new_n661_), .A3(new_n1577_), .ZN(new_n1580_));
  NAND2_X1  g1138(.A1(new_n1579_), .A2(new_n1580_), .ZN(G419));
  NAND2_X1  g1139(.A1(new_n1579_), .A2(new_n1580_), .ZN(G471));
  NAND3_X1  g1140(.A1(new_n856_), .A2(new_n861_), .A3(new_n846_), .ZN(new_n1583_));
  INV_X1    g1141(.A(new_n779_), .ZN(new_n1584_));
  AOI21_X1  g1142(.A(new_n1583_), .B1(new_n1584_), .B2(new_n1193_), .ZN(new_n1585_));
  INV_X1    g1143(.A(new_n784_), .ZN(new_n1586_));
  XNOR2_X1  g1144(.A(new_n1585_), .B(new_n1586_), .ZN(G359));
  NAND3_X1  g1145(.A1(new_n1189_), .A2(new_n1190_), .A3(new_n809_), .ZN(new_n1588_));
  AOI21_X1  g1146(.A(new_n849_), .B1(new_n1588_), .B2(new_n845_), .ZN(new_n1589_));
  INV_X1    g1147(.A(new_n1589_), .ZN(new_n1590_));
  INV_X1    g1148(.A(new_n793_), .ZN(new_n1591_));
  OAI21_X1  g1149(.A(new_n791_), .B1(new_n779_), .B2(new_n1591_), .ZN(new_n1592_));
  NAND2_X1  g1150(.A1(new_n851_), .A2(new_n810_), .ZN(new_n1593_));
  INV_X1    g1151(.A(new_n1593_), .ZN(new_n1594_));
  AOI21_X1  g1152(.A(new_n1590_), .B1(new_n1592_), .B2(new_n1594_), .ZN(new_n1595_));
  XNOR2_X1  g1153(.A(new_n1595_), .B(new_n814_), .ZN(G362));
  NAND3_X1  g1154(.A1(new_n1584_), .A2(KEYINPUT93), .A3(new_n802_), .ZN(new_n1597_));
  AOI21_X1  g1155(.A(new_n845_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n1598_));
  INV_X1    g1156(.A(KEYINPUT93), .ZN(new_n1599_));
  OAI21_X1  g1157(.A(new_n1599_), .B1(new_n779_), .B2(new_n1188_), .ZN(new_n1600_));
  NAND3_X1  g1158(.A1(new_n1597_), .A2(new_n1598_), .A3(new_n1600_), .ZN(new_n1601_));
  XNOR2_X1  g1159(.A(new_n1601_), .B(new_n1191_), .ZN(G365));
  XNOR2_X1  g1160(.A(new_n1592_), .B(new_n801_), .ZN(G368));
  NAND2_X1  g1161(.A1(new_n871_), .A2(new_n832_), .ZN(new_n1604_));
  NAND3_X1  g1162(.A1(new_n831_), .A2(new_n823_), .A3(new_n1604_), .ZN(new_n1605_));
  XNOR2_X1  g1163(.A(new_n1605_), .B(KEYINPUT94), .ZN(new_n1606_));
  NAND2_X1  g1164(.A1(new_n1606_), .A2(new_n870_), .ZN(new_n1607_));
  NOR2_X1   g1165(.A1(new_n816_), .A2(new_n865_), .ZN(new_n1608_));
  MUX2_X1   g1166(.A(new_n1607_), .B(new_n874_), .S(new_n1608_), .Z(new_n1609_));
  NAND2_X1  g1167(.A1(new_n840_), .A2(new_n841_), .ZN(new_n1610_));
  XNOR2_X1  g1168(.A(new_n1609_), .B(new_n1610_), .ZN(G347));
  OAI211_X1 g1169(.A(new_n824_), .B(new_n836_), .C1(new_n816_), .C2(new_n865_), .ZN(new_n1612_));
  INV_X1    g1170(.A(new_n872_), .ZN(new_n1613_));
  OAI211_X1 g1171(.A(new_n1612_), .B(new_n868_), .C1(new_n1185_), .C2(new_n1613_), .ZN(new_n1614_));
  XOR2_X1   g1172(.A(new_n1614_), .B(new_n831_), .Z(G350));
  NAND2_X1  g1173(.A1(new_n871_), .A2(G4420), .ZN(new_n1616_));
  INV_X1    g1174(.A(new_n1616_), .ZN(new_n1617_));
  OAI21_X1  g1175(.A(new_n1613_), .B1(new_n1608_), .B2(new_n1617_), .ZN(new_n1618_));
  XNOR2_X1  g1176(.A(new_n1618_), .B(new_n1185_), .ZN(G353));
  XNOR2_X1  g1177(.A(new_n1608_), .B(new_n836_), .ZN(G356));
  INV_X1    g1178(.A(KEYINPUT108), .ZN(new_n1621_));
  AND2_X1   g1179(.A1(new_n585_), .A2(new_n600_), .ZN(new_n1622_));
  NAND2_X1  g1180(.A1(new_n594_), .A2(new_n588_), .ZN(new_n1623_));
  NAND3_X1  g1181(.A1(new_n593_), .A2(new_n587_), .A3(new_n586_), .ZN(new_n1624_));
  AOI21_X1  g1182(.A(new_n600_), .B1(new_n1623_), .B2(new_n1624_), .ZN(new_n1625_));
  NOR2_X1   g1183(.A1(new_n1622_), .A2(new_n1625_), .ZN(new_n1626_));
  INV_X1    g1184(.A(new_n1626_), .ZN(new_n1627_));
  NAND2_X1  g1185(.A1(new_n613_), .A2(new_n1627_), .ZN(new_n1628_));
  INV_X1    g1186(.A(new_n1628_), .ZN(new_n1629_));
  NOR2_X1   g1187(.A1(new_n613_), .A2(new_n1627_), .ZN(new_n1630_));
  OAI211_X1 g1188(.A(KEYINPUT104), .B(new_n589_), .C1(new_n1629_), .C2(new_n1630_), .ZN(new_n1631_));
  NAND2_X1  g1189(.A1(new_n1543_), .A2(new_n1626_), .ZN(new_n1632_));
  INV_X1    g1190(.A(new_n589_), .ZN(new_n1633_));
  NAND3_X1  g1191(.A1(new_n1632_), .A2(new_n1633_), .A3(new_n1628_), .ZN(new_n1634_));
  NAND3_X1  g1192(.A1(new_n1631_), .A2(new_n1546_), .A3(new_n1634_), .ZN(new_n1635_));
  NAND2_X1  g1193(.A1(new_n1632_), .A2(new_n1628_), .ZN(new_n1636_));
  AOI21_X1  g1194(.A(KEYINPUT104), .B1(new_n1636_), .B2(new_n589_), .ZN(new_n1637_));
  OAI21_X1  g1195(.A(KEYINPUT105), .B1(new_n1635_), .B2(new_n1637_), .ZN(new_n1638_));
  AND2_X1   g1196(.A1(new_n1634_), .A2(new_n1546_), .ZN(new_n1639_));
  OAI21_X1  g1197(.A(new_n589_), .B1(new_n1629_), .B2(new_n1630_), .ZN(new_n1640_));
  INV_X1    g1198(.A(KEYINPUT104), .ZN(new_n1641_));
  NAND2_X1  g1199(.A1(new_n1640_), .A2(new_n1641_), .ZN(new_n1642_));
  INV_X1    g1200(.A(KEYINPUT105), .ZN(new_n1643_));
  NAND4_X1  g1201(.A1(new_n1639_), .A2(new_n1642_), .A3(new_n1643_), .A4(new_n1631_), .ZN(new_n1644_));
  AOI21_X1  g1202(.A(new_n1546_), .B1(new_n1640_), .B2(new_n1634_), .ZN(new_n1645_));
  INV_X1    g1203(.A(new_n1645_), .ZN(new_n1646_));
  NAND3_X1  g1204(.A1(new_n1638_), .A2(new_n1644_), .A3(new_n1646_), .ZN(new_n1647_));
  INV_X1    g1205(.A(KEYINPUT106), .ZN(new_n1648_));
  NAND2_X1  g1206(.A1(new_n580_), .A2(new_n1648_), .ZN(new_n1649_));
  INV_X1    g1207(.A(new_n580_), .ZN(new_n1650_));
  NAND2_X1  g1208(.A1(new_n1650_), .A2(KEYINPUT106), .ZN(new_n1651_));
  NAND3_X1  g1209(.A1(new_n1647_), .A2(new_n1649_), .A3(new_n1651_), .ZN(new_n1652_));
  NAND3_X1  g1210(.A1(new_n1639_), .A2(new_n1642_), .A3(new_n1631_), .ZN(new_n1653_));
  AOI21_X1  g1211(.A(new_n1645_), .B1(new_n1653_), .B2(KEYINPUT105), .ZN(new_n1654_));
  NAND4_X1  g1212(.A1(new_n1654_), .A2(new_n1648_), .A3(new_n580_), .A4(new_n1644_), .ZN(new_n1655_));
  INV_X1    g1213(.A(new_n572_), .ZN(new_n1656_));
  NAND4_X1  g1214(.A1(new_n1652_), .A2(new_n1655_), .A3(new_n1208_), .A4(new_n1656_), .ZN(new_n1657_));
  INV_X1    g1215(.A(KEYINPUT103), .ZN(new_n1658_));
  AOI21_X1  g1216(.A(new_n585_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n1659_));
  AOI21_X1  g1217(.A(new_n1659_), .B1(new_n585_), .B2(new_n1624_), .ZN(new_n1660_));
  AND2_X1   g1218(.A1(new_n1540_), .A2(new_n1660_), .ZN(new_n1661_));
  NOR2_X1   g1219(.A1(new_n1540_), .A2(new_n1660_), .ZN(new_n1662_));
  XNOR2_X1  g1220(.A(new_n605_), .B(new_n1561_), .ZN(new_n1663_));
  OR3_X1    g1221(.A1(new_n1661_), .A2(new_n1662_), .A3(new_n1663_), .ZN(new_n1664_));
  OAI21_X1  g1222(.A(new_n1663_), .B1(new_n1661_), .B2(new_n1662_), .ZN(new_n1665_));
  AND4_X1   g1223(.A1(KEYINPUT102), .A2(new_n1664_), .A3(new_n580_), .A4(new_n1665_), .ZN(new_n1666_));
  XOR2_X1   g1224(.A(new_n580_), .B(KEYINPUT102), .Z(new_n1667_));
  INV_X1    g1225(.A(new_n1667_), .ZN(new_n1668_));
  AOI21_X1  g1226(.A(new_n1668_), .B1(new_n1664_), .B2(new_n1665_), .ZN(new_n1669_));
  NOR3_X1   g1227(.A1(new_n1666_), .A2(new_n1669_), .A3(new_n1656_), .ZN(new_n1670_));
  NAND3_X1  g1228(.A1(new_n1208_), .A2(new_n1658_), .A3(new_n1670_), .ZN(new_n1671_));
  INV_X1    g1229(.A(new_n1671_), .ZN(new_n1672_));
  AOI21_X1  g1230(.A(new_n1658_), .B1(new_n1208_), .B2(new_n1670_), .ZN(new_n1673_));
  OAI21_X1  g1231(.A(new_n1657_), .B1(new_n1672_), .B2(new_n1673_), .ZN(new_n1674_));
  NAND2_X1  g1232(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1675_));
  INV_X1    g1233(.A(new_n1200_), .ZN(new_n1676_));
  NAND2_X1  g1234(.A1(new_n1675_), .A2(new_n1676_), .ZN(new_n1677_));
  OR2_X1    g1235(.A1(new_n1666_), .A2(new_n1669_), .ZN(new_n1678_));
  NOR2_X1   g1236(.A1(new_n572_), .A2(new_n892_), .ZN(new_n1679_));
  INV_X1    g1237(.A(new_n1679_), .ZN(new_n1680_));
  NAND2_X1  g1238(.A1(new_n1678_), .A2(new_n1680_), .ZN(new_n1681_));
  NAND2_X1  g1239(.A1(new_n1677_), .A2(new_n1681_), .ZN(new_n1682_));
  NAND2_X1  g1240(.A1(new_n1652_), .A2(new_n1655_), .ZN(new_n1683_));
  AOI21_X1  g1241(.A(new_n1682_), .B1(new_n1679_), .B2(new_n1683_), .ZN(new_n1684_));
  OAI21_X1  g1242(.A(KEYINPUT107), .B1(new_n1674_), .B2(new_n1684_), .ZN(new_n1685_));
  NAND2_X1  g1243(.A1(new_n1683_), .A2(new_n1679_), .ZN(new_n1686_));
  INV_X1    g1244(.A(new_n1682_), .ZN(new_n1687_));
  NAND2_X1  g1245(.A1(new_n1686_), .A2(new_n1687_), .ZN(new_n1688_));
  INV_X1    g1246(.A(new_n1673_), .ZN(new_n1689_));
  NAND2_X1  g1247(.A1(new_n1689_), .A2(new_n1671_), .ZN(new_n1690_));
  INV_X1    g1248(.A(KEYINPUT107), .ZN(new_n1691_));
  NAND4_X1  g1249(.A1(new_n1688_), .A2(new_n1690_), .A3(new_n1691_), .A4(new_n1657_), .ZN(new_n1692_));
  AND2_X1   g1250(.A1(new_n1685_), .A2(new_n1692_), .ZN(new_n1693_));
  NAND2_X1  g1251(.A1(new_n881_), .A2(new_n884_), .ZN(new_n1694_));
  NOR2_X1   g1252(.A1(new_n560_), .A2(new_n526_), .ZN(new_n1695_));
  NAND2_X1  g1253(.A1(new_n1291_), .A2(new_n886_), .ZN(new_n1696_));
  NAND3_X1  g1254(.A1(new_n538_), .A2(G2211), .A3(new_n539_), .ZN(new_n1697_));
  NAND3_X1  g1255(.A1(new_n1696_), .A2(new_n533_), .A3(new_n1697_), .ZN(new_n1698_));
  OAI22_X1  g1256(.A1(new_n1489_), .A2(new_n1698_), .B1(new_n544_), .B2(new_n560_), .ZN(new_n1699_));
  OAI21_X1  g1257(.A(new_n568_), .B1(new_n1489_), .B2(new_n1481_), .ZN(new_n1700_));
  NOR2_X1   g1258(.A1(new_n1699_), .A2(new_n1700_), .ZN(new_n1701_));
  AOI21_X1  g1259(.A(new_n1695_), .B1(new_n1701_), .B2(KEYINPUT95), .ZN(new_n1702_));
  INV_X1    g1260(.A(KEYINPUT95), .ZN(new_n1703_));
  OAI21_X1  g1261(.A(new_n1703_), .B1(new_n1699_), .B2(new_n1700_), .ZN(new_n1704_));
  NAND2_X1  g1262(.A1(new_n533_), .A2(new_n543_), .ZN(new_n1705_));
  AOI21_X1  g1263(.A(new_n888_), .B1(new_n531_), .B2(new_n1705_), .ZN(new_n1706_));
  AOI21_X1  g1264(.A(new_n1697_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n1707_));
  OAI211_X1 g1265(.A(new_n1698_), .B(new_n1502_), .C1(new_n1706_), .C2(new_n1707_), .ZN(new_n1708_));
  INV_X1    g1266(.A(new_n1707_), .ZN(new_n1709_));
  NAND4_X1  g1267(.A1(new_n1698_), .A2(new_n1498_), .A3(new_n1499_), .A4(new_n1500_), .ZN(new_n1710_));
  AOI21_X1  g1268(.A(new_n1492_), .B1(new_n530_), .B2(new_n528_), .ZN(new_n1711_));
  OAI211_X1 g1269(.A(new_n1709_), .B(new_n1710_), .C1(new_n1711_), .C2(new_n888_), .ZN(new_n1712_));
  AOI22_X1  g1270(.A1(new_n1702_), .A2(new_n1704_), .B1(new_n1708_), .B2(new_n1712_), .ZN(new_n1713_));
  NAND3_X1  g1271(.A1(new_n1694_), .A2(new_n1492_), .A3(new_n540_), .ZN(new_n1714_));
  NAND4_X1  g1272(.A1(new_n1483_), .A2(KEYINPUT95), .A3(new_n891_), .A4(new_n1714_), .ZN(new_n1715_));
  INV_X1    g1273(.A(new_n1695_), .ZN(new_n1716_));
  NAND3_X1  g1274(.A1(new_n1704_), .A2(new_n1715_), .A3(new_n1716_), .ZN(new_n1717_));
  NAND2_X1  g1275(.A1(new_n1708_), .A2(new_n1712_), .ZN(new_n1718_));
  NOR2_X1   g1276(.A1(new_n1717_), .A2(new_n1718_), .ZN(new_n1719_));
  OAI21_X1  g1277(.A(new_n1462_), .B1(new_n1713_), .B2(new_n1719_), .ZN(new_n1720_));
  NAND4_X1  g1278(.A1(new_n1702_), .A2(new_n1704_), .A3(new_n1708_), .A4(new_n1712_), .ZN(new_n1721_));
  NAND2_X1  g1279(.A1(new_n1717_), .A2(new_n1718_), .ZN(new_n1722_));
  NAND3_X1  g1280(.A1(new_n1721_), .A2(new_n1486_), .A3(new_n1722_), .ZN(new_n1723_));
  NAND3_X1  g1281(.A1(new_n1720_), .A2(KEYINPUT96), .A3(new_n1723_), .ZN(new_n1724_));
  INV_X1    g1282(.A(KEYINPUT96), .ZN(new_n1725_));
  NAND4_X1  g1283(.A1(new_n1721_), .A2(new_n1725_), .A3(new_n1722_), .A4(new_n1486_), .ZN(new_n1726_));
  NAND3_X1  g1284(.A1(new_n1724_), .A2(new_n533_), .A3(new_n1726_), .ZN(new_n1727_));
  NAND2_X1  g1285(.A1(new_n1727_), .A2(new_n879_), .ZN(new_n1728_));
  INV_X1    g1286(.A(KEYINPUT97), .ZN(new_n1729_));
  NAND3_X1  g1287(.A1(new_n1720_), .A2(new_n1729_), .A3(new_n1723_), .ZN(new_n1730_));
  OAI211_X1 g1288(.A(KEYINPUT97), .B(new_n1462_), .C1(new_n1713_), .C2(new_n1719_), .ZN(new_n1731_));
  AOI21_X1  g1289(.A(new_n533_), .B1(new_n1730_), .B2(new_n1731_), .ZN(new_n1732_));
  OAI21_X1  g1290(.A(new_n543_), .B1(new_n1728_), .B2(new_n1732_), .ZN(new_n1733_));
  INV_X1    g1291(.A(new_n1733_), .ZN(new_n1734_));
  INV_X1    g1292(.A(KEYINPUT98), .ZN(new_n1735_));
  NAND2_X1  g1293(.A1(new_n1724_), .A2(new_n1726_), .ZN(new_n1736_));
  NAND2_X1  g1294(.A1(new_n1736_), .A2(new_n889_), .ZN(new_n1737_));
  NAND3_X1  g1295(.A1(new_n1730_), .A2(new_n533_), .A3(new_n1731_), .ZN(new_n1738_));
  NAND2_X1  g1296(.A1(new_n1737_), .A2(new_n1738_), .ZN(new_n1739_));
  AOI21_X1  g1297(.A(new_n1735_), .B1(new_n1739_), .B2(new_n566_), .ZN(new_n1740_));
  AND3_X1   g1298(.A1(new_n1730_), .A2(new_n533_), .A3(new_n1731_), .ZN(new_n1741_));
  AOI21_X1  g1299(.A(new_n533_), .B1(new_n1724_), .B2(new_n1726_), .ZN(new_n1742_));
  OAI211_X1 g1300(.A(new_n1735_), .B(new_n566_), .C1(new_n1741_), .C2(new_n1742_), .ZN(new_n1743_));
  INV_X1    g1301(.A(new_n1743_), .ZN(new_n1744_));
  OAI21_X1  g1302(.A(new_n1734_), .B1(new_n1740_), .B2(new_n1744_), .ZN(new_n1745_));
  OAI21_X1  g1303(.A(new_n566_), .B1(new_n1741_), .B2(new_n1742_), .ZN(new_n1746_));
  NAND3_X1  g1304(.A1(new_n1737_), .A2(new_n879_), .A3(new_n1738_), .ZN(new_n1747_));
  AOI21_X1  g1305(.A(new_n543_), .B1(new_n1746_), .B2(new_n1747_), .ZN(new_n1748_));
  INV_X1    g1306(.A(new_n1748_), .ZN(new_n1749_));
  AOI21_X1  g1307(.A(new_n1694_), .B1(new_n1745_), .B2(new_n1749_), .ZN(new_n1750_));
  NAND2_X1  g1308(.A1(new_n1746_), .A2(KEYINPUT98), .ZN(new_n1751_));
  AOI21_X1  g1309(.A(new_n1733_), .B1(new_n1751_), .B2(new_n1743_), .ZN(new_n1752_));
  NOR3_X1   g1310(.A1(new_n1752_), .A2(new_n560_), .A3(new_n1748_), .ZN(new_n1753_));
  OAI21_X1  g1311(.A(new_n1677_), .B1(new_n1750_), .B2(new_n1753_), .ZN(new_n1754_));
  INV_X1    g1312(.A(KEYINPUT99), .ZN(new_n1755_));
  AOI21_X1  g1313(.A(new_n1755_), .B1(new_n531_), .B2(new_n1696_), .ZN(new_n1756_));
  OAI21_X1  g1314(.A(new_n1756_), .B1(new_n1696_), .B2(new_n1711_), .ZN(new_n1757_));
  NAND2_X1  g1315(.A1(new_n531_), .A2(new_n1705_), .ZN(new_n1758_));
  NAND3_X1  g1316(.A1(new_n1758_), .A2(new_n1755_), .A3(new_n540_), .ZN(new_n1759_));
  NAND2_X1  g1317(.A1(new_n1757_), .A2(new_n1759_), .ZN(new_n1760_));
  AOI21_X1  g1318(.A(new_n889_), .B1(new_n1485_), .B2(new_n1483_), .ZN(new_n1761_));
  NOR3_X1   g1319(.A1(new_n1700_), .A2(new_n1484_), .A3(new_n533_), .ZN(new_n1762_));
  OAI21_X1  g1320(.A(new_n1760_), .B1(new_n1761_), .B2(new_n1762_), .ZN(new_n1763_));
  NAND3_X1  g1321(.A1(new_n1485_), .A2(new_n889_), .A3(new_n1483_), .ZN(new_n1764_));
  OAI21_X1  g1322(.A(new_n533_), .B1(new_n1700_), .B2(new_n1484_), .ZN(new_n1765_));
  NAND4_X1  g1323(.A1(new_n1764_), .A2(new_n1765_), .A3(new_n1759_), .A4(new_n1757_), .ZN(new_n1766_));
  NAND3_X1  g1324(.A1(new_n1763_), .A2(new_n1486_), .A3(new_n1766_), .ZN(new_n1767_));
  INV_X1    g1325(.A(new_n1767_), .ZN(new_n1768_));
  AOI21_X1  g1326(.A(new_n1486_), .B1(new_n1763_), .B2(new_n1766_), .ZN(new_n1769_));
  NOR3_X1   g1327(.A1(new_n1768_), .A2(new_n1769_), .A3(new_n1501_), .ZN(new_n1770_));
  NAND2_X1  g1328(.A1(new_n1763_), .A2(new_n1766_), .ZN(new_n1771_));
  NAND2_X1  g1329(.A1(new_n1771_), .A2(new_n1462_), .ZN(new_n1772_));
  AOI21_X1  g1330(.A(new_n1502_), .B1(new_n1772_), .B2(new_n1767_), .ZN(new_n1773_));
  OAI21_X1  g1331(.A(new_n566_), .B1(new_n1770_), .B2(new_n1773_), .ZN(new_n1774_));
  INV_X1    g1332(.A(KEYINPUT100), .ZN(new_n1775_));
  OAI21_X1  g1333(.A(new_n1501_), .B1(new_n1768_), .B2(new_n1769_), .ZN(new_n1776_));
  NAND3_X1  g1334(.A1(new_n1772_), .A2(new_n1502_), .A3(new_n1767_), .ZN(new_n1777_));
  NAND3_X1  g1335(.A1(new_n1776_), .A2(new_n1777_), .A3(new_n879_), .ZN(new_n1778_));
  NAND3_X1  g1336(.A1(new_n1774_), .A2(new_n1775_), .A3(new_n1778_), .ZN(new_n1779_));
  NAND4_X1  g1337(.A1(new_n1776_), .A2(new_n1777_), .A3(KEYINPUT100), .A4(new_n879_), .ZN(new_n1780_));
  NAND3_X1  g1338(.A1(new_n1779_), .A2(new_n880_), .A3(new_n1780_), .ZN(new_n1781_));
  NAND4_X1  g1339(.A1(new_n1774_), .A2(KEYINPUT101), .A3(new_n543_), .A4(new_n1778_), .ZN(new_n1782_));
  NAND3_X1  g1340(.A1(new_n1774_), .A2(new_n543_), .A3(new_n1778_), .ZN(new_n1783_));
  INV_X1    g1341(.A(KEYINPUT101), .ZN(new_n1784_));
  NAND2_X1  g1342(.A1(new_n1783_), .A2(new_n1784_), .ZN(new_n1785_));
  NAND3_X1  g1343(.A1(new_n1781_), .A2(new_n1782_), .A3(new_n1785_), .ZN(new_n1786_));
  NAND2_X1  g1344(.A1(new_n1786_), .A2(new_n560_), .ZN(new_n1787_));
  NAND4_X1  g1345(.A1(new_n1781_), .A2(new_n1785_), .A3(new_n1694_), .A4(new_n1782_), .ZN(new_n1788_));
  NAND3_X1  g1346(.A1(new_n1787_), .A2(new_n1208_), .A3(new_n1788_), .ZN(new_n1789_));
  AOI21_X1  g1347(.A(new_n1693_), .B1(new_n1754_), .B2(new_n1789_), .ZN(new_n1790_));
  NAND3_X1  g1348(.A1(new_n1688_), .A2(new_n1690_), .A3(new_n1657_), .ZN(new_n1791_));
  NAND2_X1  g1349(.A1(new_n1789_), .A2(new_n1791_), .ZN(new_n1792_));
  NAND3_X1  g1350(.A1(new_n1745_), .A2(new_n1694_), .A3(new_n1749_), .ZN(new_n1793_));
  NAND2_X1  g1351(.A1(new_n1746_), .A2(new_n1747_), .ZN(new_n1794_));
  AOI21_X1  g1352(.A(new_n1694_), .B1(new_n1794_), .B2(new_n543_), .ZN(new_n1795_));
  NOR2_X1   g1353(.A1(new_n1740_), .A2(new_n1744_), .ZN(new_n1796_));
  OAI21_X1  g1354(.A(new_n880_), .B1(new_n1728_), .B2(new_n1732_), .ZN(new_n1797_));
  OAI21_X1  g1355(.A(new_n1795_), .B1(new_n1796_), .B2(new_n1797_), .ZN(new_n1798_));
  NAND2_X1  g1356(.A1(new_n1793_), .A2(new_n1798_), .ZN(new_n1799_));
  AOI21_X1  g1357(.A(new_n1792_), .B1(new_n1677_), .B2(new_n1799_), .ZN(new_n1800_));
  OAI21_X1  g1358(.A(new_n1621_), .B1(new_n1790_), .B2(new_n1800_), .ZN(new_n1801_));
  NAND2_X1  g1359(.A1(new_n1799_), .A2(new_n1677_), .ZN(new_n1802_));
  AND2_X1   g1360(.A1(new_n1789_), .A2(new_n1791_), .ZN(new_n1803_));
  NAND2_X1  g1361(.A1(new_n1802_), .A2(new_n1803_), .ZN(new_n1804_));
  OAI21_X1  g1362(.A(new_n560_), .B1(new_n1752_), .B2(new_n1748_), .ZN(new_n1805_));
  AOI21_X1  g1363(.A(new_n1208_), .B1(new_n1793_), .B2(new_n1805_), .ZN(new_n1806_));
  INV_X1    g1364(.A(new_n1789_), .ZN(new_n1807_));
  NOR2_X1   g1365(.A1(new_n1806_), .A2(new_n1807_), .ZN(new_n1808_));
  OAI211_X1 g1366(.A(new_n1804_), .B(KEYINPUT108), .C1(new_n1808_), .C2(new_n1693_), .ZN(new_n1809_));
  NAND2_X1  g1367(.A1(new_n1801_), .A2(new_n1809_), .ZN(G321));
  OAI21_X1  g1368(.A(new_n680_), .B1(new_n676_), .B2(new_n631_), .ZN(new_n1811_));
  NAND2_X1  g1369(.A1(new_n1811_), .A2(new_n636_), .ZN(new_n1812_));
  AOI21_X1  g1370(.A(new_n1515_), .B1(new_n675_), .B2(new_n1517_), .ZN(new_n1813_));
  NAND3_X1  g1371(.A1(new_n1813_), .A2(new_n637_), .A3(new_n1519_), .ZN(new_n1814_));
  NAND2_X1  g1372(.A1(new_n1812_), .A2(new_n1814_), .ZN(new_n1815_));
  INV_X1    g1373(.A(KEYINPUT109), .ZN(new_n1816_));
  NAND3_X1  g1374(.A1(new_n672_), .A2(new_n676_), .A3(new_n1816_), .ZN(new_n1817_));
  OAI21_X1  g1375(.A(KEYINPUT109), .B1(new_n671_), .B2(new_n675_), .ZN(new_n1818_));
  AOI21_X1  g1376(.A(new_n646_), .B1(new_n1817_), .B2(new_n1818_), .ZN(new_n1819_));
  OR2_X1    g1377(.A1(new_n1815_), .A2(new_n1819_), .ZN(new_n1820_));
  NAND2_X1  g1378(.A1(new_n1511_), .A2(new_n647_), .ZN(new_n1821_));
  INV_X1    g1379(.A(new_n1821_), .ZN(new_n1822_));
  NAND2_X1  g1380(.A1(new_n1815_), .A2(new_n1819_), .ZN(new_n1823_));
  AND3_X1   g1381(.A1(new_n1820_), .A2(new_n1822_), .A3(new_n1823_), .ZN(new_n1824_));
  AND2_X1   g1382(.A1(new_n1812_), .A2(new_n1814_), .ZN(new_n1825_));
  NAND2_X1  g1383(.A1(new_n1819_), .A2(KEYINPUT110), .ZN(new_n1826_));
  NAND2_X1  g1384(.A1(new_n1825_), .A2(new_n1826_), .ZN(new_n1827_));
  NAND3_X1  g1385(.A1(new_n1815_), .A2(new_n1819_), .A3(KEYINPUT110), .ZN(new_n1828_));
  AOI21_X1  g1386(.A(new_n1822_), .B1(new_n1827_), .B2(new_n1828_), .ZN(new_n1829_));
  NOR3_X1   g1387(.A1(new_n1824_), .A2(new_n1829_), .A3(new_n639_), .ZN(new_n1830_));
  NAND2_X1  g1388(.A1(new_n1827_), .A2(new_n1828_), .ZN(new_n1831_));
  NAND2_X1  g1389(.A1(new_n1831_), .A2(new_n1821_), .ZN(new_n1832_));
  NAND3_X1  g1390(.A1(new_n1820_), .A2(new_n1822_), .A3(new_n1823_), .ZN(new_n1833_));
  AOI21_X1  g1391(.A(new_n1467_), .B1(new_n1832_), .B2(new_n1833_), .ZN(new_n1834_));
  OAI21_X1  g1392(.A(new_n645_), .B1(new_n1830_), .B2(new_n1834_), .ZN(new_n1835_));
  NAND3_X1  g1393(.A1(new_n1832_), .A2(new_n1467_), .A3(new_n1833_), .ZN(new_n1836_));
  NAND2_X1  g1394(.A1(new_n1831_), .A2(new_n1822_), .ZN(new_n1837_));
  NAND3_X1  g1395(.A1(new_n1820_), .A2(new_n1821_), .A3(new_n1823_), .ZN(new_n1838_));
  NAND3_X1  g1396(.A1(new_n1837_), .A2(new_n639_), .A3(new_n1838_), .ZN(new_n1839_));
  NAND3_X1  g1397(.A1(new_n1836_), .A2(new_n1839_), .A3(new_n1518_), .ZN(new_n1840_));
  NAND3_X1  g1398(.A1(new_n1835_), .A2(new_n655_), .A3(new_n1840_), .ZN(new_n1841_));
  INV_X1    g1399(.A(new_n1841_), .ZN(new_n1842_));
  AOI21_X1  g1400(.A(new_n655_), .B1(new_n1835_), .B2(new_n1840_), .ZN(new_n1843_));
  OAI21_X1  g1401(.A(new_n631_), .B1(new_n1842_), .B2(new_n1843_), .ZN(new_n1844_));
  NAND2_X1  g1402(.A1(new_n1844_), .A2(KEYINPUT111), .ZN(new_n1845_));
  NAND2_X1  g1403(.A1(new_n1835_), .A2(new_n1840_), .ZN(new_n1846_));
  NAND2_X1  g1404(.A1(new_n1846_), .A2(new_n656_), .ZN(new_n1847_));
  NAND2_X1  g1405(.A1(new_n1847_), .A2(new_n1841_), .ZN(new_n1848_));
  INV_X1    g1406(.A(KEYINPUT111), .ZN(new_n1849_));
  NAND3_X1  g1407(.A1(new_n1848_), .A2(new_n1849_), .A3(new_n631_), .ZN(new_n1850_));
  NAND2_X1  g1408(.A1(new_n1845_), .A2(new_n1850_), .ZN(new_n1851_));
  OAI21_X1  g1409(.A(new_n1518_), .B1(new_n1830_), .B2(new_n1834_), .ZN(new_n1852_));
  NAND3_X1  g1410(.A1(new_n1836_), .A2(new_n1839_), .A3(new_n645_), .ZN(new_n1853_));
  NAND3_X1  g1411(.A1(new_n1852_), .A2(new_n656_), .A3(new_n1853_), .ZN(new_n1854_));
  NAND3_X1  g1412(.A1(new_n1841_), .A2(new_n1854_), .A3(new_n1517_), .ZN(new_n1855_));
  XNOR2_X1  g1413(.A(new_n1855_), .B(KEYINPUT112), .ZN(new_n1856_));
  NAND3_X1  g1414(.A1(new_n1851_), .A2(new_n678_), .A3(new_n1856_), .ZN(new_n1857_));
  NAND2_X1  g1415(.A1(new_n1848_), .A2(new_n1517_), .ZN(new_n1858_));
  NAND3_X1  g1416(.A1(new_n1841_), .A2(new_n1854_), .A3(new_n631_), .ZN(new_n1859_));
  NAND3_X1  g1417(.A1(new_n1858_), .A2(new_n623_), .A3(new_n1859_), .ZN(new_n1860_));
  AOI21_X1  g1418(.A(new_n1475_), .B1(new_n1857_), .B2(new_n1860_), .ZN(new_n1861_));
  AND2_X1   g1419(.A1(new_n1813_), .A2(new_n638_), .ZN(new_n1862_));
  AOI21_X1  g1420(.A(new_n1509_), .B1(new_n1813_), .B2(new_n1519_), .ZN(new_n1863_));
  NOR2_X1   g1421(.A1(new_n1862_), .A2(new_n1863_), .ZN(new_n1864_));
  NAND2_X1  g1422(.A1(new_n1817_), .A2(new_n1818_), .ZN(new_n1865_));
  NOR2_X1   g1423(.A1(new_n1864_), .A2(new_n1865_), .ZN(new_n1866_));
  INV_X1    g1424(.A(new_n1865_), .ZN(new_n1867_));
  NOR3_X1   g1425(.A1(new_n1867_), .A2(new_n1862_), .A3(new_n1863_), .ZN(new_n1868_));
  OAI21_X1  g1426(.A(new_n1512_), .B1(new_n1866_), .B2(new_n1868_), .ZN(new_n1869_));
  NAND2_X1  g1427(.A1(new_n1864_), .A2(new_n1865_), .ZN(new_n1870_));
  OAI21_X1  g1428(.A(new_n643_), .B1(new_n1509_), .B2(new_n645_), .ZN(new_n1871_));
  OAI21_X1  g1429(.A(new_n1871_), .B1(new_n1862_), .B2(new_n1863_), .ZN(new_n1872_));
  NAND3_X1  g1430(.A1(new_n1870_), .A2(new_n1511_), .A3(new_n1872_), .ZN(new_n1873_));
  NAND3_X1  g1431(.A1(new_n1869_), .A2(new_n1467_), .A3(new_n1873_), .ZN(new_n1874_));
  INV_X1    g1432(.A(new_n1874_), .ZN(new_n1875_));
  AOI21_X1  g1433(.A(new_n1467_), .B1(new_n1869_), .B2(new_n1873_), .ZN(new_n1876_));
  OAI21_X1  g1434(.A(new_n1518_), .B1(new_n1875_), .B2(new_n1876_), .ZN(new_n1877_));
  OAI21_X1  g1435(.A(new_n1511_), .B1(new_n1866_), .B2(new_n1868_), .ZN(new_n1878_));
  NAND3_X1  g1436(.A1(new_n1870_), .A2(new_n1512_), .A3(new_n1872_), .ZN(new_n1879_));
  NAND3_X1  g1437(.A1(new_n1878_), .A2(new_n639_), .A3(new_n1879_), .ZN(new_n1880_));
  NAND3_X1  g1438(.A1(new_n1874_), .A2(new_n1880_), .A3(new_n645_), .ZN(new_n1881_));
  AND4_X1   g1439(.A1(new_n656_), .A2(new_n1877_), .A3(new_n1517_), .A4(new_n1881_), .ZN(new_n1882_));
  OAI21_X1  g1440(.A(new_n645_), .B1(new_n1875_), .B2(new_n1876_), .ZN(new_n1883_));
  NAND3_X1  g1441(.A1(new_n1874_), .A2(new_n1880_), .A3(new_n1518_), .ZN(new_n1884_));
  NAND3_X1  g1442(.A1(new_n1883_), .A2(new_n655_), .A3(new_n1884_), .ZN(new_n1885_));
  AOI21_X1  g1443(.A(new_n655_), .B1(new_n1883_), .B2(new_n1884_), .ZN(new_n1886_));
  NAND2_X1  g1444(.A1(new_n631_), .A2(KEYINPUT113), .ZN(new_n1887_));
  OAI21_X1  g1445(.A(new_n1885_), .B1(new_n1886_), .B2(new_n1887_), .ZN(new_n1888_));
  INV_X1    g1446(.A(new_n1887_), .ZN(new_n1889_));
  NAND4_X1  g1447(.A1(new_n1883_), .A2(new_n1884_), .A3(new_n655_), .A4(new_n1889_), .ZN(new_n1890_));
  AOI21_X1  g1448(.A(new_n1882_), .B1(new_n1888_), .B2(new_n1890_), .ZN(new_n1891_));
  NOR2_X1   g1449(.A1(new_n1891_), .A2(new_n678_), .ZN(new_n1892_));
  AOI211_X1 g1450(.A(new_n623_), .B(new_n1882_), .C1(new_n1888_), .C2(new_n1890_), .ZN(new_n1893_));
  OAI21_X1  g1451(.A(new_n1475_), .B1(new_n1892_), .B2(new_n1893_), .ZN(new_n1894_));
  AND2_X1   g1452(.A1(new_n685_), .A2(new_n1569_), .ZN(new_n1895_));
  NAND2_X1  g1453(.A1(new_n1475_), .A2(new_n1895_), .ZN(new_n1896_));
  XNOR2_X1  g1454(.A(new_n1896_), .B(KEYINPUT114), .ZN(new_n1897_));
  NAND2_X1  g1455(.A1(new_n685_), .A2(new_n658_), .ZN(new_n1898_));
  AOI22_X1  g1456(.A1(new_n1895_), .A2(new_n658_), .B1(new_n1898_), .B2(new_n1572_), .ZN(new_n1899_));
  NAND2_X1  g1457(.A1(new_n684_), .A2(new_n1572_), .ZN(new_n1900_));
  MUX2_X1   g1458(.A(new_n1899_), .B(new_n1900_), .S(new_n1475_), .Z(new_n1901_));
  NAND2_X1  g1459(.A1(new_n1897_), .A2(new_n1901_), .ZN(new_n1902_));
  NAND2_X1  g1460(.A1(new_n1894_), .A2(new_n1902_), .ZN(new_n1903_));
  NOR2_X1   g1461(.A1(new_n1861_), .A2(new_n1903_), .ZN(new_n1904_));
  AND3_X1   g1462(.A1(new_n1851_), .A2(new_n678_), .A3(new_n1856_), .ZN(new_n1905_));
  AOI21_X1  g1463(.A(new_n678_), .B1(new_n1851_), .B2(new_n1856_), .ZN(new_n1906_));
  OAI21_X1  g1464(.A(new_n1476_), .B1(new_n1905_), .B2(new_n1906_), .ZN(new_n1907_));
  NAND2_X1  g1465(.A1(new_n1907_), .A2(new_n1894_), .ZN(new_n1908_));
  INV_X1    g1466(.A(new_n1902_), .ZN(new_n1909_));
  AOI21_X1  g1467(.A(new_n1904_), .B1(new_n1908_), .B2(new_n1909_), .ZN(G338));
  NAND4_X1  g1468(.A1(new_n856_), .A2(new_n861_), .A3(new_n815_), .A4(new_n846_), .ZN(new_n1911_));
  NAND2_X1  g1469(.A1(new_n1590_), .A2(new_n1591_), .ZN(new_n1912_));
  NAND2_X1  g1470(.A1(new_n1598_), .A2(new_n1188_), .ZN(new_n1913_));
  NAND3_X1  g1471(.A1(new_n1589_), .A2(new_n793_), .A3(new_n1593_), .ZN(new_n1914_));
  NAND3_X1  g1472(.A1(new_n1912_), .A2(new_n1913_), .A3(new_n1914_), .ZN(new_n1915_));
  INV_X1    g1473(.A(new_n1915_), .ZN(new_n1916_));
  AOI21_X1  g1474(.A(new_n1913_), .B1(new_n1912_), .B2(new_n1914_), .ZN(new_n1917_));
  OAI21_X1  g1475(.A(new_n1911_), .B1(new_n1916_), .B2(new_n1917_), .ZN(new_n1918_));
  INV_X1    g1476(.A(new_n1917_), .ZN(new_n1919_));
  NAND2_X1  g1477(.A1(new_n1919_), .A2(new_n1915_), .ZN(new_n1920_));
  XNOR2_X1  g1478(.A(new_n1911_), .B(KEYINPUT115), .ZN(new_n1921_));
  OAI211_X1 g1479(.A(new_n1918_), .B(new_n1563_), .C1(new_n1920_), .C2(new_n1921_), .ZN(new_n1922_));
  NAND3_X1  g1480(.A1(new_n1919_), .A2(new_n1915_), .A3(new_n1911_), .ZN(new_n1923_));
  NOR2_X1   g1481(.A1(new_n1916_), .A2(new_n1917_), .ZN(new_n1924_));
  OAI211_X1 g1482(.A(new_n1923_), .B(new_n794_), .C1(new_n1924_), .C2(new_n1921_), .ZN(new_n1925_));
  NAND2_X1  g1483(.A1(new_n1922_), .A2(new_n1925_), .ZN(new_n1926_));
  NAND2_X1  g1484(.A1(new_n1926_), .A2(new_n851_), .ZN(new_n1927_));
  OAI21_X1  g1485(.A(new_n1918_), .B1(new_n1920_), .B2(new_n1921_), .ZN(new_n1928_));
  NAND2_X1  g1486(.A1(new_n1928_), .A2(new_n794_), .ZN(new_n1929_));
  NAND3_X1  g1487(.A1(new_n1929_), .A2(new_n801_), .A3(new_n1922_), .ZN(new_n1930_));
  AOI21_X1  g1488(.A(new_n784_), .B1(new_n1927_), .B2(new_n1930_), .ZN(new_n1931_));
  INV_X1    g1489(.A(new_n1931_), .ZN(new_n1932_));
  NAND2_X1  g1490(.A1(new_n1929_), .A2(new_n1922_), .ZN(new_n1933_));
  NAND2_X1  g1491(.A1(new_n1933_), .A2(new_n851_), .ZN(new_n1934_));
  INV_X1    g1492(.A(KEYINPUT116), .ZN(new_n1935_));
  NAND3_X1  g1493(.A1(new_n1922_), .A2(new_n1925_), .A3(new_n801_), .ZN(new_n1936_));
  NAND4_X1  g1494(.A1(new_n1934_), .A2(new_n1935_), .A3(new_n862_), .A4(new_n1936_), .ZN(new_n1937_));
  NAND2_X1  g1495(.A1(new_n1936_), .A2(new_n862_), .ZN(new_n1938_));
  AOI21_X1  g1496(.A(new_n801_), .B1(new_n1929_), .B2(new_n1922_), .ZN(new_n1939_));
  OAI21_X1  g1497(.A(KEYINPUT116), .B1(new_n1938_), .B2(new_n1939_), .ZN(new_n1940_));
  NAND4_X1  g1498(.A1(new_n1932_), .A2(new_n1937_), .A3(new_n810_), .A4(new_n1940_), .ZN(new_n1941_));
  AND3_X1   g1499(.A1(new_n1927_), .A2(new_n1930_), .A3(new_n784_), .ZN(new_n1942_));
  OAI21_X1  g1500(.A(new_n1191_), .B1(new_n1942_), .B2(new_n1931_), .ZN(new_n1943_));
  NAND3_X1  g1501(.A1(new_n1941_), .A2(new_n814_), .A3(new_n1943_), .ZN(new_n1944_));
  NOR3_X1   g1502(.A1(new_n1942_), .A2(new_n1931_), .A3(new_n1191_), .ZN(new_n1945_));
  NAND3_X1  g1503(.A1(new_n1932_), .A2(new_n1937_), .A3(new_n1940_), .ZN(new_n1946_));
  AOI21_X1  g1504(.A(new_n1945_), .B1(new_n854_), .B2(new_n1946_), .ZN(new_n1947_));
  OAI21_X1  g1505(.A(new_n1944_), .B1(new_n1947_), .B2(new_n814_), .ZN(new_n1948_));
  AOI21_X1  g1506(.A(new_n778_), .B1(new_n741_), .B2(new_n1187_), .ZN(new_n1949_));
  INV_X1    g1507(.A(new_n1949_), .ZN(new_n1950_));
  NAND2_X1  g1508(.A1(new_n1948_), .A2(new_n1950_), .ZN(new_n1951_));
  INV_X1    g1509(.A(KEYINPUT118), .ZN(new_n1952_));
  NAND2_X1  g1510(.A1(new_n1912_), .A2(new_n791_), .ZN(new_n1953_));
  AOI21_X1  g1511(.A(new_n1953_), .B1(new_n793_), .B2(new_n1589_), .ZN(new_n1954_));
  OR2_X1    g1512(.A1(new_n1598_), .A2(new_n1191_), .ZN(new_n1955_));
  AOI21_X1  g1513(.A(new_n791_), .B1(new_n1955_), .B2(new_n850_), .ZN(new_n1956_));
  OR2_X1    g1514(.A1(new_n1954_), .A2(new_n1956_), .ZN(new_n1957_));
  NAND2_X1  g1515(.A1(new_n856_), .A2(new_n861_), .ZN(new_n1958_));
  NAND2_X1  g1516(.A1(new_n1958_), .A2(new_n1598_), .ZN(new_n1959_));
  OAI21_X1  g1517(.A(new_n1959_), .B1(new_n1583_), .B2(new_n1598_), .ZN(new_n1960_));
  NAND2_X1  g1518(.A1(new_n1960_), .A2(new_n851_), .ZN(new_n1961_));
  INV_X1    g1519(.A(new_n1961_), .ZN(new_n1962_));
  NOR2_X1   g1520(.A1(new_n1960_), .A2(new_n851_), .ZN(new_n1963_));
  OAI21_X1  g1521(.A(new_n1957_), .B1(new_n1962_), .B2(new_n1963_), .ZN(new_n1964_));
  INV_X1    g1522(.A(new_n1963_), .ZN(new_n1965_));
  NOR2_X1   g1523(.A1(new_n1954_), .A2(new_n1956_), .ZN(new_n1966_));
  NAND3_X1  g1524(.A1(new_n1965_), .A2(new_n1961_), .A3(new_n1966_), .ZN(new_n1967_));
  AND3_X1   g1525(.A1(new_n1964_), .A2(new_n1586_), .A3(new_n1967_), .ZN(new_n1968_));
  AOI21_X1  g1526(.A(new_n1194_), .B1(new_n1964_), .B2(new_n1967_), .ZN(new_n1969_));
  OR3_X1    g1527(.A1(new_n1968_), .A2(new_n1969_), .A3(new_n854_), .ZN(new_n1970_));
  AOI21_X1  g1528(.A(new_n1586_), .B1(new_n1964_), .B2(new_n1967_), .ZN(new_n1971_));
  OAI21_X1  g1529(.A(new_n1191_), .B1(new_n1968_), .B2(new_n1971_), .ZN(new_n1972_));
  NAND2_X1  g1530(.A1(new_n1970_), .A2(new_n1972_), .ZN(new_n1973_));
  NAND2_X1  g1531(.A1(new_n1973_), .A2(new_n1192_), .ZN(new_n1974_));
  NAND3_X1  g1532(.A1(new_n1970_), .A2(new_n814_), .A3(new_n1972_), .ZN(new_n1975_));
  NAND3_X1  g1533(.A1(new_n1974_), .A2(new_n1949_), .A3(new_n1975_), .ZN(new_n1976_));
  XOR2_X1   g1534(.A(new_n1610_), .B(new_n836_), .Z(new_n1977_));
  XNOR2_X1  g1535(.A(new_n1977_), .B(new_n874_), .ZN(new_n1978_));
  MUX2_X1   g1536(.A(new_n821_), .B(new_n822_), .S(new_n872_), .Z(new_n1979_));
  XNOR2_X1  g1537(.A(new_n1978_), .B(new_n1979_), .ZN(new_n1980_));
  NOR2_X1   g1538(.A1(new_n1980_), .A2(new_n824_), .ZN(new_n1981_));
  AOI21_X1  g1539(.A(new_n1981_), .B1(new_n823_), .B2(new_n1980_), .ZN(new_n1982_));
  OR2_X1    g1540(.A1(new_n1982_), .A2(new_n831_), .ZN(new_n1983_));
  NAND2_X1  g1541(.A1(new_n1982_), .A2(new_n831_), .ZN(new_n1984_));
  XOR2_X1   g1542(.A(new_n864_), .B(KEYINPUT117), .Z(new_n1985_));
  OAI21_X1  g1543(.A(new_n1950_), .B1(new_n1985_), .B2(new_n1201_), .ZN(new_n1986_));
  NAND2_X1  g1544(.A1(new_n1949_), .A2(new_n1985_), .ZN(new_n1987_));
  NAND4_X1  g1545(.A1(new_n1983_), .A2(new_n1984_), .A3(new_n1986_), .A4(new_n1987_), .ZN(new_n1988_));
  AOI22_X1  g1546(.A1(new_n1617_), .A2(new_n821_), .B1(new_n822_), .B2(new_n1604_), .ZN(new_n1989_));
  XNOR2_X1  g1547(.A(new_n1977_), .B(new_n1989_), .ZN(new_n1990_));
  XNOR2_X1  g1548(.A(new_n1990_), .B(new_n1607_), .ZN(new_n1991_));
  NAND2_X1  g1549(.A1(new_n1991_), .A2(new_n823_), .ZN(new_n1992_));
  OAI21_X1  g1550(.A(new_n1992_), .B1(new_n824_), .B2(new_n1991_), .ZN(new_n1993_));
  XNOR2_X1  g1551(.A(new_n1993_), .B(new_n831_), .ZN(new_n1994_));
  OAI21_X1  g1552(.A(new_n1986_), .B1(new_n864_), .B2(new_n1950_), .ZN(new_n1995_));
  NAND2_X1  g1553(.A1(new_n1994_), .A2(new_n1995_), .ZN(new_n1996_));
  NAND2_X1  g1554(.A1(new_n1988_), .A2(new_n1996_), .ZN(new_n1997_));
  AND2_X1   g1555(.A1(new_n1976_), .A2(new_n1997_), .ZN(new_n1998_));
  AND3_X1   g1556(.A1(new_n1951_), .A2(new_n1952_), .A3(new_n1998_), .ZN(new_n1999_));
  AOI21_X1  g1557(.A(new_n1952_), .B1(new_n1951_), .B2(new_n1998_), .ZN(new_n2000_));
  INV_X1    g1558(.A(new_n1944_), .ZN(new_n2001_));
  AOI21_X1  g1559(.A(new_n814_), .B1(new_n1941_), .B2(new_n1943_), .ZN(new_n2002_));
  OAI21_X1  g1560(.A(new_n1950_), .B1(new_n2001_), .B2(new_n2002_), .ZN(new_n2003_));
  AOI21_X1  g1561(.A(new_n1997_), .B1(new_n2003_), .B2(new_n1976_), .ZN(new_n2004_));
  NOR3_X1   g1562(.A1(new_n1999_), .A2(new_n2000_), .A3(new_n2004_), .ZN(G370));
  AND2_X1   g1563(.A1(new_n719_), .A2(new_n723_), .ZN(new_n2006_));
  NAND2_X1  g1564(.A1(new_n2006_), .A2(new_n738_), .ZN(new_n2007_));
  NAND3_X1  g1565(.A1(new_n709_), .A2(new_n1238_), .A3(new_n730_), .ZN(new_n2008_));
  NAND2_X1  g1566(.A1(new_n2007_), .A2(new_n2008_), .ZN(new_n2009_));
  OAI211_X1 g1567(.A(new_n2009_), .B(new_n697_), .C1(new_n725_), .C2(new_n731_), .ZN(new_n2010_));
  NAND2_X1  g1568(.A1(new_n732_), .A2(new_n2007_), .ZN(new_n2011_));
  NAND2_X1  g1569(.A1(new_n1222_), .A2(new_n503_), .ZN(new_n2012_));
  INV_X1    g1570(.A(new_n503_), .ZN(new_n2013_));
  NAND2_X1  g1571(.A1(new_n1224_), .A2(new_n2013_), .ZN(new_n2014_));
  OAI21_X1  g1572(.A(new_n2012_), .B1(new_n2014_), .B2(new_n1222_), .ZN(new_n2015_));
  AND3_X1   g1573(.A1(new_n2010_), .A2(new_n2011_), .A3(new_n2015_), .ZN(new_n2016_));
  AOI21_X1  g1574(.A(new_n2015_), .B1(new_n2010_), .B2(new_n2011_), .ZN(new_n2017_));
  OAI21_X1  g1575(.A(new_n1210_), .B1(new_n2016_), .B2(new_n2017_), .ZN(new_n2018_));
  NAND2_X1  g1576(.A1(new_n2010_), .A2(new_n2011_), .ZN(new_n2019_));
  INV_X1    g1577(.A(new_n2015_), .ZN(new_n2020_));
  NAND2_X1  g1578(.A1(new_n2019_), .A2(new_n2020_), .ZN(new_n2021_));
  NAND3_X1  g1579(.A1(new_n2010_), .A2(new_n2011_), .A3(new_n2015_), .ZN(new_n2022_));
  NAND3_X1  g1580(.A1(new_n2021_), .A2(new_n2022_), .A3(new_n504_), .ZN(new_n2023_));
  NAND3_X1  g1581(.A1(new_n2018_), .A2(new_n2023_), .A3(KEYINPUT119), .ZN(new_n2024_));
  INV_X1    g1582(.A(KEYINPUT119), .ZN(new_n2025_));
  OAI211_X1 g1583(.A(new_n2025_), .B(new_n1210_), .C1(new_n2016_), .C2(new_n2017_), .ZN(new_n2026_));
  NAND3_X1  g1584(.A1(new_n2024_), .A2(new_n1211_), .A3(new_n2026_), .ZN(new_n2027_));
  AND2_X1   g1585(.A1(new_n2018_), .A2(new_n2023_), .ZN(new_n2028_));
  NAND2_X1  g1586(.A1(new_n2028_), .A2(new_n1223_), .ZN(new_n2029_));
  AND3_X1   g1587(.A1(new_n2027_), .A2(new_n2029_), .A3(new_n1217_), .ZN(new_n2030_));
  AOI21_X1  g1588(.A(new_n1217_), .B1(new_n2027_), .B2(new_n2029_), .ZN(new_n2031_));
  OAI21_X1  g1589(.A(new_n705_), .B1(new_n2030_), .B2(new_n2031_), .ZN(new_n2032_));
  NAND3_X1  g1590(.A1(new_n2027_), .A2(new_n2029_), .A3(new_n1217_), .ZN(new_n2033_));
  NAND3_X1  g1591(.A1(new_n2024_), .A2(new_n1223_), .A3(new_n2026_), .ZN(new_n2034_));
  NAND2_X1  g1592(.A1(new_n2028_), .A2(new_n1211_), .ZN(new_n2035_));
  NAND3_X1  g1593(.A1(new_n2034_), .A2(new_n2035_), .A3(new_n737_), .ZN(new_n2036_));
  NAND3_X1  g1594(.A1(new_n2033_), .A2(new_n2036_), .A3(new_n709_), .ZN(new_n2037_));
  NAND3_X1  g1595(.A1(new_n2032_), .A2(new_n730_), .A3(new_n2037_), .ZN(new_n2038_));
  INV_X1    g1596(.A(new_n2038_), .ZN(new_n2039_));
  AOI21_X1  g1597(.A(new_n730_), .B1(new_n2032_), .B2(new_n2037_), .ZN(new_n2040_));
  OAI21_X1  g1598(.A(G4526), .B1(new_n2039_), .B2(new_n2040_), .ZN(new_n2041_));
  NAND2_X1  g1599(.A1(new_n2041_), .A2(KEYINPUT127), .ZN(new_n2042_));
  INV_X1    g1600(.A(KEYINPUT127), .ZN(new_n2043_));
  OAI211_X1 g1601(.A(new_n2043_), .B(G4526), .C1(new_n2039_), .C2(new_n2040_), .ZN(new_n2044_));
  INV_X1    g1602(.A(new_n705_), .ZN(new_n2045_));
  NAND2_X1  g1603(.A1(new_n1222_), .A2(new_n501_), .ZN(new_n2046_));
  OAI211_X1 g1604(.A(new_n1221_), .B(new_n1226_), .C1(new_n723_), .C2(new_n705_), .ZN(new_n2047_));
  NAND3_X1  g1605(.A1(new_n1232_), .A2(new_n1235_), .A3(new_n2045_), .ZN(new_n2048_));
  NAND3_X1  g1606(.A1(new_n2046_), .A2(new_n2047_), .A3(new_n2048_), .ZN(new_n2049_));
  AND2_X1   g1607(.A1(new_n2049_), .A2(new_n724_), .ZN(new_n2050_));
  NOR2_X1   g1608(.A1(new_n2049_), .A2(new_n724_), .ZN(new_n2051_));
  OAI21_X1  g1609(.A(new_n732_), .B1(new_n2050_), .B2(new_n2051_), .ZN(new_n2052_));
  INV_X1    g1610(.A(KEYINPUT120), .ZN(new_n2053_));
  NAND2_X1  g1611(.A1(new_n2052_), .A2(new_n2053_), .ZN(new_n2054_));
  OAI211_X1 g1612(.A(KEYINPUT120), .B(new_n732_), .C1(new_n2050_), .C2(new_n2051_), .ZN(new_n2055_));
  NAND2_X1  g1613(.A1(new_n2054_), .A2(new_n2055_), .ZN(new_n2056_));
  NOR2_X1   g1614(.A1(new_n2050_), .A2(new_n2051_), .ZN(new_n2057_));
  INV_X1    g1615(.A(KEYINPUT121), .ZN(new_n2058_));
  NAND2_X1  g1616(.A1(new_n732_), .A2(new_n2058_), .ZN(new_n2059_));
  OAI211_X1 g1617(.A(KEYINPUT121), .B(new_n697_), .C1(new_n725_), .C2(new_n731_), .ZN(new_n2060_));
  NAND2_X1  g1618(.A1(new_n2059_), .A2(new_n2060_), .ZN(new_n2061_));
  AND3_X1   g1619(.A1(new_n2057_), .A2(KEYINPUT122), .A3(new_n2061_), .ZN(new_n2062_));
  AOI21_X1  g1620(.A(KEYINPUT122), .B1(new_n2057_), .B2(new_n2061_), .ZN(new_n2063_));
  OAI21_X1  g1621(.A(new_n2056_), .B1(new_n2062_), .B2(new_n2063_), .ZN(new_n2064_));
  NAND2_X1  g1622(.A1(new_n2064_), .A2(new_n1210_), .ZN(new_n2065_));
  OAI211_X1 g1623(.A(new_n2056_), .B(new_n504_), .C1(new_n2063_), .C2(new_n2062_), .ZN(new_n2066_));
  AOI21_X1  g1624(.A(new_n1223_), .B1(new_n2065_), .B2(new_n2066_), .ZN(new_n2067_));
  OAI21_X1  g1625(.A(KEYINPUT123), .B1(new_n2057_), .B2(new_n2061_), .ZN(new_n2068_));
  NAND2_X1  g1626(.A1(new_n2057_), .A2(new_n1215_), .ZN(new_n2069_));
  NAND2_X1  g1627(.A1(new_n2068_), .A2(new_n2069_), .ZN(new_n2070_));
  NOR3_X1   g1628(.A1(new_n2057_), .A2(new_n2061_), .A3(KEYINPUT123), .ZN(new_n2071_));
  OAI21_X1  g1629(.A(new_n1210_), .B1(new_n2070_), .B2(new_n2071_), .ZN(new_n2072_));
  AND3_X1   g1630(.A1(new_n2072_), .A2(new_n2066_), .A3(new_n1223_), .ZN(new_n2073_));
  OAI21_X1  g1631(.A(new_n737_), .B1(new_n2067_), .B2(new_n2073_), .ZN(new_n2074_));
  INV_X1    g1632(.A(new_n2066_), .ZN(new_n2075_));
  NAND2_X1  g1633(.A1(new_n2057_), .A2(new_n2061_), .ZN(new_n2076_));
  INV_X1    g1634(.A(KEYINPUT122), .ZN(new_n2077_));
  NAND2_X1  g1635(.A1(new_n2076_), .A2(new_n2077_), .ZN(new_n2078_));
  NAND3_X1  g1636(.A1(new_n2057_), .A2(KEYINPUT122), .A3(new_n2061_), .ZN(new_n2079_));
  NAND2_X1  g1637(.A1(new_n2078_), .A2(new_n2079_), .ZN(new_n2080_));
  AOI21_X1  g1638(.A(new_n504_), .B1(new_n2080_), .B2(new_n2056_), .ZN(new_n2081_));
  OAI21_X1  g1639(.A(new_n1211_), .B1(new_n2075_), .B2(new_n2081_), .ZN(new_n2082_));
  NAND3_X1  g1640(.A1(new_n2072_), .A2(new_n2066_), .A3(new_n1223_), .ZN(new_n2083_));
  NAND3_X1  g1641(.A1(new_n2082_), .A2(new_n1217_), .A3(new_n2083_), .ZN(new_n2084_));
  AOI21_X1  g1642(.A(new_n2045_), .B1(new_n2074_), .B2(new_n2084_), .ZN(new_n2085_));
  INV_X1    g1643(.A(KEYINPUT124), .ZN(new_n2086_));
  NOR3_X1   g1644(.A1(new_n2067_), .A2(new_n2073_), .A3(new_n737_), .ZN(new_n2087_));
  NAND3_X1  g1645(.A1(new_n2072_), .A2(new_n2066_), .A3(new_n1211_), .ZN(new_n2088_));
  NAND2_X1  g1646(.A1(new_n2088_), .A2(new_n737_), .ZN(new_n2089_));
  AOI21_X1  g1647(.A(new_n1211_), .B1(new_n2065_), .B2(new_n2066_), .ZN(new_n2090_));
  OAI21_X1  g1648(.A(new_n709_), .B1(new_n2089_), .B2(new_n2090_), .ZN(new_n2091_));
  OAI21_X1  g1649(.A(new_n2086_), .B1(new_n2087_), .B2(new_n2091_), .ZN(new_n2092_));
  OAI21_X1  g1650(.A(new_n1223_), .B1(new_n2075_), .B2(new_n2081_), .ZN(new_n2093_));
  NAND3_X1  g1651(.A1(new_n2093_), .A2(new_n737_), .A3(new_n2088_), .ZN(new_n2094_));
  NAND4_X1  g1652(.A1(new_n2084_), .A2(new_n2094_), .A3(KEYINPUT124), .A4(new_n709_), .ZN(new_n2095_));
  AOI21_X1  g1653(.A(new_n2085_), .B1(new_n2092_), .B2(new_n2095_), .ZN(new_n2096_));
  OAI21_X1  g1654(.A(new_n505_), .B1(new_n2096_), .B2(new_n730_), .ZN(new_n2097_));
  AOI211_X1 g1655(.A(new_n731_), .B(new_n2085_), .C1(new_n2092_), .C2(new_n2095_), .ZN(new_n2098_));
  OAI211_X1 g1656(.A(new_n2042_), .B(new_n2044_), .C1(new_n2097_), .C2(new_n2098_), .ZN(new_n2099_));
  XNOR2_X1  g1657(.A(new_n1248_), .B(new_n1254_), .ZN(new_n2100_));
  NAND2_X1  g1658(.A1(new_n770_), .A2(new_n752_), .ZN(new_n2101_));
  OAI21_X1  g1659(.A(new_n2101_), .B1(new_n760_), .B2(new_n752_), .ZN(new_n2102_));
  XOR2_X1   g1660(.A(new_n2102_), .B(new_n755_), .Z(new_n2103_));
  XNOR2_X1  g1661(.A(new_n2100_), .B(new_n2103_), .ZN(new_n2104_));
  NOR2_X1   g1662(.A1(new_n2104_), .A2(new_n1260_), .ZN(new_n2105_));
  NAND2_X1  g1663(.A1(new_n2104_), .A2(new_n1260_), .ZN(new_n2106_));
  AOI21_X1  g1664(.A(new_n2105_), .B1(KEYINPUT125), .B2(new_n2106_), .ZN(new_n2107_));
  OAI21_X1  g1665(.A(new_n2107_), .B1(KEYINPUT125), .B2(new_n2106_), .ZN(new_n2108_));
  NOR2_X1   g1666(.A1(new_n734_), .A2(G4526), .ZN(new_n2109_));
  NAND4_X1  g1667(.A1(new_n1257_), .A2(new_n773_), .A3(new_n746_), .A4(new_n747_), .ZN(new_n2110_));
  OAI21_X1  g1668(.A(new_n2110_), .B1(new_n1260_), .B2(new_n774_), .ZN(new_n2111_));
  NAND2_X1  g1669(.A1(new_n753_), .A2(new_n759_), .ZN(new_n2112_));
  AOI21_X1  g1670(.A(new_n754_), .B1(new_n2112_), .B2(new_n2101_), .ZN(new_n2113_));
  NOR2_X1   g1671(.A1(new_n2113_), .A2(new_n1256_), .ZN(new_n2114_));
  XNOR2_X1  g1672(.A(new_n2111_), .B(new_n2114_), .ZN(new_n2115_));
  XOR2_X1   g1673(.A(new_n761_), .B(new_n1254_), .Z(new_n2116_));
  XNOR2_X1  g1674(.A(new_n2115_), .B(new_n2116_), .ZN(new_n2117_));
  AOI22_X1  g1675(.A1(new_n2108_), .A2(new_n2109_), .B1(new_n742_), .B2(new_n2117_), .ZN(new_n2118_));
  OAI21_X1  g1676(.A(new_n734_), .B1(new_n737_), .B2(new_n2008_), .ZN(new_n2119_));
  INV_X1    g1677(.A(KEYINPUT126), .ZN(new_n2120_));
  OR2_X1    g1678(.A1(new_n2119_), .A2(new_n2120_), .ZN(new_n2121_));
  NAND2_X1  g1679(.A1(new_n2119_), .A2(new_n2120_), .ZN(new_n2122_));
  NAND4_X1  g1680(.A1(new_n2108_), .A2(G4526), .A3(new_n2121_), .A4(new_n2122_), .ZN(new_n2123_));
  AND2_X1   g1681(.A1(new_n2118_), .A2(new_n2123_), .ZN(new_n2124_));
  AND2_X1   g1682(.A1(new_n2092_), .A2(new_n2095_), .ZN(new_n2125_));
  OAI21_X1  g1683(.A(new_n731_), .B1(new_n2125_), .B2(new_n2085_), .ZN(new_n2126_));
  NAND2_X1  g1684(.A1(new_n2096_), .A2(new_n730_), .ZN(new_n2127_));
  NAND3_X1  g1685(.A1(new_n2126_), .A2(new_n505_), .A3(new_n2127_), .ZN(new_n2128_));
  NOR3_X1   g1686(.A1(new_n2030_), .A2(new_n2031_), .A3(new_n705_), .ZN(new_n2129_));
  AOI21_X1  g1687(.A(new_n709_), .B1(new_n2036_), .B2(new_n2033_), .ZN(new_n2130_));
  OAI21_X1  g1688(.A(new_n731_), .B1(new_n2129_), .B2(new_n2130_), .ZN(new_n2131_));
  NAND2_X1  g1689(.A1(new_n2131_), .A2(new_n2038_), .ZN(new_n2132_));
  AOI21_X1  g1690(.A(new_n2124_), .B1(new_n2132_), .B2(G4526), .ZN(new_n2133_));
  AOI22_X1  g1691(.A1(new_n2099_), .A2(new_n2124_), .B1(new_n2128_), .B2(new_n2133_), .ZN(G399));
endmodule


