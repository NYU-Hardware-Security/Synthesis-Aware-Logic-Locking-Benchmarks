//Secret key is'1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_c6288" written by ABC on Sun Nov 20 20:03:01 2022

module locked_c6288 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G18gat, G35gat,
    G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat,
    G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat,
    G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat,
    G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat,
    G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat,
    G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat,
    G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_n129_, new_n130_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_;
  INV_X1    g0000(.A(G1gat), .ZN(new_n129_));
  INV_X1    g0001(.A(G273gat), .ZN(new_n130_));
  NOR2_X1   g0002(.A1(new_n129_), .A2(new_n130_), .ZN(G545gat));
  INV_X1    g0003(.A(G18gat), .ZN(new_n132_));
  INV_X1    g0004(.A(G290gat), .ZN(new_n133_));
  NOR4_X1   g0005(.A1(new_n129_), .A2(new_n132_), .A3(new_n130_), .A4(new_n133_), .ZN(new_n134_));
  AOI22_X1  g0006(.A1(G1gat), .A2(G290gat), .B1(G18gat), .B2(G273gat), .ZN(new_n135_));
  NOR2_X1   g0007(.A1(new_n134_), .A2(new_n135_), .ZN(G1581gat));
  NAND4_X1  g0008(.A1(G18gat), .A2(G35gat), .A3(G273gat), .A4(G290gat), .ZN(new_n137_));
  AOI22_X1  g0009(.A1(G18gat), .A2(G290gat), .B1(G35gat), .B2(G273gat), .ZN(new_n138_));
  OAI21_X1  g0010(.A(new_n137_), .B1(new_n138_), .B2(KEYINPUT0), .ZN(new_n139_));
  AOI21_X1  g0011(.A(new_n139_), .B1(KEYINPUT0), .B2(new_n138_), .ZN(new_n140_));
  XOR2_X1   g0012(.A(new_n140_), .B(new_n134_), .Z(new_n141_));
  NAND2_X1  g0013(.A1(G1gat), .A2(G307gat), .ZN(new_n142_));
  XNOR2_X1  g0014(.A(new_n141_), .B(new_n142_), .ZN(G1901gat));
  NAND2_X1  g0015(.A1(new_n141_), .A2(new_n142_), .ZN(new_n144_));
  NAND4_X1  g0016(.A1(G35gat), .A2(G52gat), .A3(G273gat), .A4(G290gat), .ZN(new_n145_));
  INV_X1    g0017(.A(new_n145_), .ZN(new_n146_));
  AOI22_X1  g0018(.A1(G35gat), .A2(G290gat), .B1(G52gat), .B2(G273gat), .ZN(new_n147_));
  OAI21_X1  g0019(.A(new_n137_), .B1(new_n146_), .B2(new_n147_), .ZN(new_n148_));
  OAI21_X1  g0020(.A(new_n148_), .B1(new_n137_), .B2(new_n146_), .ZN(new_n149_));
  INV_X1    g0021(.A(G307gat), .ZN(new_n150_));
  NOR2_X1   g0022(.A1(new_n132_), .A2(new_n150_), .ZN(new_n151_));
  XOR2_X1   g0023(.A(new_n149_), .B(new_n151_), .Z(new_n152_));
  INV_X1    g0024(.A(new_n152_), .ZN(new_n153_));
  OR2_X1    g0025(.A1(new_n140_), .A2(new_n134_), .ZN(new_n154_));
  NAND3_X1  g0026(.A1(new_n144_), .A2(new_n153_), .A3(new_n154_), .ZN(new_n155_));
  INV_X1    g0027(.A(new_n155_), .ZN(new_n156_));
  AOI21_X1  g0028(.A(new_n153_), .B1(new_n144_), .B2(new_n154_), .ZN(new_n157_));
  NOR2_X1   g0029(.A1(new_n156_), .A2(new_n157_), .ZN(new_n158_));
  INV_X1    g0030(.A(G324gat), .ZN(new_n159_));
  NOR2_X1   g0031(.A1(new_n129_), .A2(new_n159_), .ZN(new_n160_));
  INV_X1    g0032(.A(new_n160_), .ZN(new_n161_));
  XNOR2_X1  g0033(.A(new_n158_), .B(new_n161_), .ZN(G2223gat));
  AOI21_X1  g0034(.A(new_n157_), .B1(new_n161_), .B2(new_n155_), .ZN(new_n163_));
  INV_X1    g0035(.A(new_n163_), .ZN(new_n164_));
  INV_X1    g0036(.A(G52gat), .ZN(new_n165_));
  INV_X1    g0037(.A(G69gat), .ZN(new_n166_));
  OAI22_X1  g0038(.A1(new_n165_), .A2(new_n133_), .B1(new_n166_), .B2(new_n130_), .ZN(new_n167_));
  NAND4_X1  g0039(.A1(G52gat), .A2(G69gat), .A3(G273gat), .A4(G290gat), .ZN(new_n168_));
  AOI21_X1  g0040(.A(new_n146_), .B1(new_n167_), .B2(new_n168_), .ZN(new_n169_));
  AOI21_X1  g0041(.A(new_n169_), .B1(new_n146_), .B2(new_n168_), .ZN(new_n170_));
  NAND2_X1  g0042(.A1(G35gat), .A2(G307gat), .ZN(new_n171_));
  OR2_X1    g0043(.A1(new_n170_), .A2(new_n171_), .ZN(new_n172_));
  NAND2_X1  g0044(.A1(new_n170_), .A2(new_n171_), .ZN(new_n173_));
  NAND2_X1  g0045(.A1(new_n172_), .A2(new_n173_), .ZN(new_n174_));
  NOR2_X1   g0046(.A1(new_n146_), .A2(new_n137_), .ZN(new_n175_));
  OAI21_X1  g0047(.A(new_n148_), .B1(new_n175_), .B2(new_n151_), .ZN(new_n176_));
  INV_X1    g0048(.A(new_n176_), .ZN(new_n177_));
  NOR2_X1   g0049(.A1(new_n174_), .A2(new_n177_), .ZN(new_n178_));
  INV_X1    g0050(.A(new_n178_), .ZN(new_n179_));
  NOR2_X1   g0051(.A1(new_n132_), .A2(new_n159_), .ZN(new_n180_));
  INV_X1    g0052(.A(new_n180_), .ZN(new_n181_));
  NAND2_X1  g0053(.A1(new_n174_), .A2(new_n177_), .ZN(new_n182_));
  NAND3_X1  g0054(.A1(new_n179_), .A2(new_n181_), .A3(new_n182_), .ZN(new_n183_));
  INV_X1    g0055(.A(new_n182_), .ZN(new_n184_));
  OAI21_X1  g0056(.A(new_n180_), .B1(new_n184_), .B2(new_n178_), .ZN(new_n185_));
  NAND3_X1  g0057(.A1(new_n164_), .A2(new_n183_), .A3(new_n185_), .ZN(new_n186_));
  NAND2_X1  g0058(.A1(new_n185_), .A2(new_n183_), .ZN(new_n187_));
  NAND2_X1  g0059(.A1(new_n187_), .A2(new_n163_), .ZN(new_n188_));
  NAND2_X1  g0060(.A1(new_n186_), .A2(new_n188_), .ZN(new_n189_));
  NAND2_X1  g0061(.A1(G1gat), .A2(G341gat), .ZN(new_n190_));
  NOR2_X1   g0062(.A1(new_n189_), .A2(new_n190_), .ZN(new_n191_));
  NAND3_X1  g0063(.A1(new_n186_), .A2(new_n190_), .A3(new_n188_), .ZN(new_n192_));
  INV_X1    g0064(.A(KEYINPUT1), .ZN(new_n193_));
  NAND2_X1  g0065(.A1(new_n192_), .A2(new_n193_), .ZN(new_n194_));
  NAND4_X1  g0066(.A1(new_n186_), .A2(KEYINPUT1), .A3(new_n190_), .A4(new_n188_), .ZN(new_n195_));
  NAND2_X1  g0067(.A1(new_n194_), .A2(new_n195_), .ZN(new_n196_));
  AOI21_X1  g0068(.A(new_n191_), .B1(new_n196_), .B2(new_n190_), .ZN(G2548gat));
  INV_X1    g0069(.A(G341gat), .ZN(new_n198_));
  NOR2_X1   g0070(.A1(new_n132_), .A2(new_n198_), .ZN(new_n199_));
  INV_X1    g0071(.A(new_n199_), .ZN(new_n200_));
  NAND2_X1  g0072(.A1(new_n183_), .A2(new_n179_), .ZN(new_n201_));
  INV_X1    g0073(.A(new_n169_), .ZN(new_n202_));
  AOI22_X1  g0074(.A1(new_n170_), .A2(new_n171_), .B1(KEYINPUT2), .B2(new_n202_), .ZN(new_n203_));
  OR2_X1    g0075(.A1(new_n202_), .A2(KEYINPUT2), .ZN(new_n204_));
  NAND2_X1  g0076(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND4_X1  g0077(.A1(G69gat), .A2(G86gat), .A3(G273gat), .A4(G290gat), .ZN(new_n206_));
  INV_X1    g0078(.A(new_n206_), .ZN(new_n207_));
  OR2_X1    g0079(.A1(new_n207_), .A2(new_n168_), .ZN(new_n208_));
  AOI22_X1  g0080(.A1(G69gat), .A2(G290gat), .B1(G86gat), .B2(G273gat), .ZN(new_n209_));
  OAI21_X1  g0081(.A(new_n168_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g0082(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g0083(.A1(new_n165_), .A2(new_n150_), .ZN(new_n212_));
  NAND2_X1  g0084(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g0085(.A(new_n212_), .ZN(new_n214_));
  NAND3_X1  g0086(.A1(new_n208_), .A2(new_n214_), .A3(new_n210_), .ZN(new_n215_));
  AND2_X1   g0087(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g0088(.A1(new_n205_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g0089(.A(G35gat), .ZN(new_n218_));
  NOR2_X1   g0090(.A1(new_n218_), .A2(new_n159_), .ZN(new_n219_));
  INV_X1    g0091(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g0092(.A1(new_n205_), .A2(new_n216_), .ZN(new_n221_));
  NAND3_X1  g0093(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g0094(.A(new_n220_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n223_));
  INV_X1    g0095(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g0096(.A(new_n201_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g0097(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g0098(.A1(new_n201_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n227_));
  AOI21_X1  g0099(.A(new_n200_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g0100(.A(new_n227_), .ZN(new_n229_));
  NOR3_X1   g0101(.A1(new_n229_), .A2(new_n225_), .A3(new_n199_), .ZN(new_n230_));
  OAI211_X1 g0102(.A(new_n186_), .B(new_n192_), .C1(new_n228_), .C2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g0103(.A1(new_n228_), .A2(new_n230_), .ZN(new_n232_));
  INV_X1    g0104(.A(new_n232_), .ZN(new_n233_));
  INV_X1    g0105(.A(new_n186_), .ZN(new_n234_));
  AOI21_X1  g0106(.A(new_n234_), .B1(new_n194_), .B2(new_n195_), .ZN(new_n235_));
  OAI21_X1  g0107(.A(new_n231_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g0108(.A1(G1gat), .A2(G358gat), .ZN(new_n237_));
  XOR2_X1   g0109(.A(new_n236_), .B(new_n237_), .Z(G2877gat));
  OAI21_X1  g0110(.A(new_n227_), .B1(new_n225_), .B2(new_n199_), .ZN(new_n239_));
  INV_X1    g0111(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g0112(.A1(new_n222_), .A2(new_n221_), .ZN(new_n241_));
  INV_X1    g0113(.A(G86gat), .ZN(new_n242_));
  INV_X1    g0114(.A(G103gat), .ZN(new_n243_));
  OAI22_X1  g0115(.A1(new_n242_), .A2(new_n133_), .B1(new_n243_), .B2(new_n130_), .ZN(new_n244_));
  NAND4_X1  g0116(.A1(G86gat), .A2(G103gat), .A3(G273gat), .A4(G290gat), .ZN(new_n245_));
  NAND2_X1  g0117(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g0118(.A1(new_n246_), .A2(new_n206_), .ZN(new_n247_));
  NAND2_X1  g0119(.A1(new_n207_), .A2(new_n245_), .ZN(new_n248_));
  NAND2_X1  g0120(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g0121(.A1(new_n166_), .A2(new_n150_), .ZN(new_n250_));
  NAND2_X1  g0122(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g0123(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g0124(.A1(new_n247_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g0125(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g0126(.A1(new_n254_), .A2(new_n210_), .A3(new_n215_), .ZN(new_n255_));
  NAND2_X1  g0127(.A1(new_n215_), .A2(new_n210_), .ZN(new_n256_));
  NAND3_X1  g0128(.A1(new_n251_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g0129(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g0130(.A1(new_n165_), .A2(new_n159_), .ZN(new_n259_));
  INV_X1    g0131(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g0132(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g0133(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n262_));
  NAND3_X1  g0134(.A1(new_n241_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g0135(.A1(new_n261_), .A2(KEYINPUT3), .A3(new_n262_), .ZN(new_n264_));
  INV_X1    g0136(.A(KEYINPUT3), .ZN(new_n265_));
  NAND3_X1  g0137(.A1(new_n258_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n266_));
  NAND4_X1  g0138(.A1(new_n264_), .A2(new_n221_), .A3(new_n222_), .A4(new_n266_), .ZN(new_n267_));
  NOR2_X1   g0139(.A1(new_n218_), .A2(new_n198_), .ZN(new_n268_));
  NAND3_X1  g0140(.A1(new_n263_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g0141(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g0142(.A(new_n268_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n271_));
  OAI21_X1  g0143(.A(new_n240_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g0144(.A(new_n271_), .ZN(new_n273_));
  NAND3_X1  g0145(.A1(new_n239_), .A2(new_n273_), .A3(new_n269_), .ZN(new_n274_));
  NAND2_X1  g0146(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g0147(.A(G358gat), .ZN(new_n276_));
  NOR2_X1   g0148(.A1(new_n132_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g0149(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g0150(.A(new_n275_), .B(new_n278_), .ZN(new_n279_));
  OAI211_X1 g0151(.A(new_n237_), .B(new_n231_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n280_));
  INV_X1    g0152(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g0153(.A(KEYINPUT4), .ZN(new_n282_));
  NOR2_X1   g0154(.A1(new_n235_), .A2(new_n282_), .ZN(new_n283_));
  AOI211_X1 g0155(.A(KEYINPUT4), .B(new_n234_), .C1(new_n194_), .C2(new_n195_), .ZN(new_n284_));
  NOR3_X1   g0156(.A1(new_n283_), .A2(new_n284_), .A3(new_n233_), .ZN(new_n285_));
  OR3_X1    g0157(.A1(new_n279_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g0158(.A(new_n279_), .B1(new_n285_), .B2(new_n281_), .ZN(new_n287_));
  NAND2_X1  g0159(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g0160(.A(G375gat), .ZN(new_n289_));
  NOR2_X1   g0161(.A1(new_n129_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g0162(.A(new_n288_), .B(new_n290_), .ZN(G3211gat));
  NOR2_X1   g0163(.A1(new_n132_), .A2(new_n289_), .ZN(new_n292_));
  INV_X1    g0164(.A(new_n272_), .ZN(new_n293_));
  OAI21_X1  g0165(.A(new_n274_), .B1(new_n293_), .B2(new_n277_), .ZN(new_n294_));
  NAND2_X1  g0166(.A1(new_n257_), .A2(new_n259_), .ZN(new_n295_));
  NAND2_X1  g0167(.A1(new_n295_), .A2(new_n255_), .ZN(new_n296_));
  INV_X1    g0168(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g0169(.A1(new_n166_), .A2(new_n159_), .ZN(new_n298_));
  INV_X1    g0170(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g0171(.A(G120gat), .ZN(new_n300_));
  OAI22_X1  g0172(.A1(new_n243_), .A2(new_n133_), .B1(new_n300_), .B2(new_n130_), .ZN(new_n301_));
  NAND4_X1  g0173(.A1(G103gat), .A2(G120gat), .A3(G273gat), .A4(G290gat), .ZN(new_n302_));
  NAND2_X1  g0174(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g0175(.A1(new_n303_), .A2(new_n245_), .ZN(new_n304_));
  NOR2_X1   g0176(.A1(new_n242_), .A2(new_n150_), .ZN(new_n305_));
  INV_X1    g0177(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g0178(.A(new_n302_), .ZN(new_n307_));
  OR2_X1    g0179(.A1(new_n307_), .A2(new_n245_), .ZN(new_n308_));
  NAND3_X1  g0180(.A1(new_n304_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g0181(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g0182(.A(new_n306_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n311_));
  OAI211_X1 g0183(.A(new_n247_), .B(new_n253_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g0184(.A1(new_n253_), .A2(new_n247_), .ZN(new_n313_));
  INV_X1    g0185(.A(new_n311_), .ZN(new_n314_));
  NAND3_X1  g0186(.A1(new_n313_), .A2(new_n314_), .A3(new_n309_), .ZN(new_n315_));
  AOI21_X1  g0187(.A(new_n299_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g0188(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g0189(.A1(new_n312_), .A2(new_n315_), .A3(new_n299_), .ZN(new_n318_));
  NAND3_X1  g0190(.A1(new_n297_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g0191(.A(new_n318_), .ZN(new_n320_));
  OAI21_X1  g0192(.A(new_n296_), .B1(new_n320_), .B2(new_n316_), .ZN(new_n321_));
  NAND2_X1  g0193(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g0194(.A1(new_n165_), .A2(new_n198_), .ZN(new_n323_));
  XOR2_X1   g0195(.A(new_n323_), .B(KEYINPUT6), .Z(new_n324_));
  OR2_X1    g0196(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g0197(.A1(new_n322_), .A2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g0198(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g0199(.A1(new_n241_), .A2(new_n266_), .A3(new_n264_), .ZN(new_n328_));
  NAND3_X1  g0200(.A1(new_n273_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  OR2_X1    g0201(.A1(new_n322_), .A2(new_n323_), .ZN(new_n330_));
  INV_X1    g0202(.A(new_n328_), .ZN(new_n331_));
  OAI211_X1 g0203(.A(new_n326_), .B(new_n330_), .C1(new_n271_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g0204(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g0205(.A1(new_n333_), .A2(G35gat), .A3(G358gat), .ZN(new_n334_));
  NAND2_X1  g0206(.A1(G35gat), .A2(G358gat), .ZN(new_n335_));
  NAND3_X1  g0207(.A1(new_n329_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  AND2_X1   g0208(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g0209(.A1(new_n274_), .A2(KEYINPUT5), .ZN(new_n338_));
  AOI21_X1  g0210(.A(new_n294_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AND4_X1   g0211(.A1(new_n294_), .A2(new_n334_), .A3(new_n338_), .A4(new_n336_), .ZN(new_n340_));
  OAI21_X1  g0212(.A(new_n292_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g0213(.A1(new_n334_), .A2(new_n338_), .A3(new_n336_), .ZN(new_n342_));
  OAI211_X1 g0214(.A(new_n342_), .B(new_n274_), .C1(new_n277_), .C2(new_n275_), .ZN(new_n343_));
  NAND3_X1  g0215(.A1(new_n337_), .A2(new_n294_), .A3(new_n338_), .ZN(new_n344_));
  INV_X1    g0216(.A(new_n292_), .ZN(new_n345_));
  NAND3_X1  g0217(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g0218(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  NOR3_X1   g0219(.A1(new_n279_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n348_));
  OAI21_X1  g0220(.A(new_n287_), .B1(new_n348_), .B2(new_n290_), .ZN(new_n349_));
  NAND2_X1  g0221(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g0222(.A1(new_n350_), .A2(KEYINPUT8), .ZN(new_n351_));
  INV_X1    g0223(.A(KEYINPUT8), .ZN(new_n352_));
  NAND3_X1  g0224(.A1(new_n347_), .A2(new_n352_), .A3(new_n349_), .ZN(new_n353_));
  NAND2_X1  g0225(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g0226(.A(new_n287_), .ZN(new_n355_));
  INV_X1    g0227(.A(new_n290_), .ZN(new_n356_));
  AOI21_X1  g0228(.A(new_n355_), .B1(new_n356_), .B2(new_n286_), .ZN(new_n357_));
  NAND4_X1  g0229(.A1(new_n357_), .A2(KEYINPUT7), .A3(new_n346_), .A4(new_n341_), .ZN(new_n358_));
  INV_X1    g0230(.A(KEYINPUT7), .ZN(new_n359_));
  OAI21_X1  g0231(.A(new_n359_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n360_));
  NAND2_X1  g0232(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g0233(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g0234(.A(G392gat), .ZN(new_n363_));
  NOR2_X1   g0235(.A1(new_n129_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g0236(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g0237(.A(new_n362_), .B(new_n365_), .ZN(G3552gat));
  NAND2_X1  g0238(.A1(new_n362_), .A2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g0239(.A1(new_n357_), .A2(new_n347_), .ZN(new_n368_));
  INV_X1    g0240(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g0241(.A1(new_n337_), .A2(new_n294_), .ZN(new_n370_));
  NAND2_X1  g0242(.A1(new_n346_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g0243(.A1(new_n370_), .A2(KEYINPUT9), .ZN(new_n372_));
  OR3_X1    g0244(.A1(new_n271_), .A2(KEYINPUT10), .A3(new_n331_), .ZN(new_n373_));
  OAI21_X1  g0245(.A(KEYINPUT10), .B1(new_n271_), .B2(new_n331_), .ZN(new_n374_));
  NAND2_X1  g0246(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g0247(.A(new_n336_), .B1(new_n375_), .B2(new_n327_), .ZN(new_n376_));
  INV_X1    g0248(.A(G137gat), .ZN(new_n377_));
  OAI22_X1  g0249(.A1(new_n300_), .A2(new_n133_), .B1(new_n377_), .B2(new_n130_), .ZN(new_n378_));
  NAND4_X1  g0250(.A1(G120gat), .A2(G137gat), .A3(G273gat), .A4(G290gat), .ZN(new_n379_));
  NAND2_X1  g0251(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g0252(.A1(new_n380_), .A2(new_n302_), .ZN(new_n381_));
  INV_X1    g0253(.A(new_n379_), .ZN(new_n382_));
  NOR2_X1   g0254(.A1(new_n382_), .A2(new_n302_), .ZN(new_n383_));
  INV_X1    g0255(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g0256(.A1(new_n243_), .A2(new_n150_), .ZN(new_n385_));
  NAND3_X1  g0257(.A1(new_n381_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g0258(.A(KEYINPUT11), .ZN(new_n387_));
  NAND2_X1  g0259(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g0260(.A(new_n385_), .ZN(new_n389_));
  INV_X1    g0261(.A(new_n381_), .ZN(new_n390_));
  OAI21_X1  g0262(.A(new_n389_), .B1(new_n390_), .B2(new_n383_), .ZN(new_n391_));
  NAND4_X1  g0263(.A1(new_n381_), .A2(new_n384_), .A3(KEYINPUT11), .A4(new_n385_), .ZN(new_n392_));
  NAND3_X1  g0264(.A1(new_n388_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AOI22_X1  g0265(.A1(new_n308_), .A2(new_n306_), .B1(new_n303_), .B2(new_n245_), .ZN(new_n394_));
  INV_X1    g0266(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g0267(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g0268(.A1(new_n242_), .A2(new_n159_), .ZN(new_n397_));
  INV_X1    g0269(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g0270(.A1(new_n391_), .A2(new_n394_), .A3(new_n386_), .ZN(new_n399_));
  NAND3_X1  g0271(.A1(new_n396_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g0272(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g0273(.A(new_n398_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n402_));
  OAI211_X1 g0274(.A(new_n315_), .B(new_n318_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  INV_X1    g0275(.A(new_n402_), .ZN(new_n404_));
  NAND2_X1  g0276(.A1(new_n318_), .A2(new_n315_), .ZN(new_n405_));
  NAND3_X1  g0277(.A1(new_n404_), .A2(new_n405_), .A3(new_n400_), .ZN(new_n406_));
  NAND2_X1  g0278(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g0279(.A1(new_n166_), .A2(new_n198_), .ZN(new_n408_));
  NAND2_X1  g0280(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g0281(.A(new_n408_), .ZN(new_n410_));
  NAND3_X1  g0282(.A1(new_n403_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n411_));
  NAND4_X1  g0283(.A1(new_n409_), .A2(new_n325_), .A3(new_n319_), .A4(new_n411_), .ZN(new_n412_));
  OAI21_X1  g0284(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n413_));
  AND3_X1   g0285(.A1(new_n403_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n414_));
  AOI21_X1  g0286(.A(new_n410_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n415_));
  OAI21_X1  g0287(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g0288(.A1(new_n165_), .A2(new_n276_), .ZN(new_n417_));
  AND3_X1   g0289(.A1(new_n412_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g0290(.A(new_n417_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n419_));
  NOR2_X1   g0291(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g0292(.A1(new_n376_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g0293(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g0294(.A1(new_n218_), .A2(new_n289_), .ZN(new_n423_));
  INV_X1    g0295(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g0296(.A1(new_n376_), .A2(new_n420_), .ZN(new_n425_));
  NAND3_X1  g0297(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g0298(.A(new_n425_), .ZN(new_n427_));
  OAI21_X1  g0299(.A(new_n423_), .B1(new_n427_), .B2(new_n421_), .ZN(new_n428_));
  NAND4_X1  g0300(.A1(new_n371_), .A2(new_n372_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n429_));
  NOR2_X1   g0301(.A1(new_n132_), .A2(new_n363_), .ZN(new_n430_));
  INV_X1    g0302(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g0303(.A1(new_n428_), .A2(new_n426_), .A3(new_n372_), .ZN(new_n432_));
  NAND3_X1  g0304(.A1(new_n432_), .A2(new_n346_), .A3(new_n370_), .ZN(new_n433_));
  NAND3_X1  g0305(.A1(new_n429_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g0306(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g0307(.A(new_n431_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n436_));
  OR2_X1    g0308(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g0309(.A1(new_n367_), .A2(new_n369_), .A3(new_n437_), .ZN(new_n438_));
  NOR2_X1   g0310(.A1(new_n435_), .A2(new_n436_), .ZN(new_n439_));
  AOI21_X1  g0311(.A(new_n364_), .B1(new_n354_), .B2(new_n361_), .ZN(new_n440_));
  OAI21_X1  g0312(.A(new_n439_), .B1(new_n440_), .B2(new_n368_), .ZN(new_n441_));
  NAND2_X1  g0313(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g0314(.A(G409gat), .ZN(new_n443_));
  NOR2_X1   g0315(.A1(new_n129_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g0316(.A(new_n442_), .B(new_n444_), .ZN(G3895gat));
  AOI21_X1  g0317(.A(new_n437_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n446_));
  INV_X1    g0318(.A(new_n444_), .ZN(new_n447_));
  AOI21_X1  g0319(.A(new_n446_), .B1(new_n447_), .B2(new_n438_), .ZN(new_n448_));
  NAND3_X1  g0320(.A1(new_n371_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n449_));
  NAND2_X1  g0321(.A1(new_n434_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g0322(.A1(new_n218_), .A2(new_n363_), .ZN(new_n451_));
  INV_X1    g0323(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g0324(.A(new_n425_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n453_));
  NOR2_X1   g0325(.A1(new_n165_), .A2(new_n289_), .ZN(new_n454_));
  INV_X1    g0326(.A(new_n454_), .ZN(new_n455_));
  AND3_X1   g0327(.A1(new_n409_), .A2(new_n413_), .A3(new_n411_), .ZN(new_n456_));
  NOR2_X1   g0328(.A1(new_n419_), .A2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g0329(.A1(new_n393_), .A2(new_n395_), .B1(new_n399_), .B2(new_n398_), .ZN(new_n458_));
  NOR2_X1   g0330(.A1(new_n243_), .A2(new_n159_), .ZN(new_n459_));
  INV_X1    g0331(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g0332(.A(new_n381_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n461_));
  NAND4_X1  g0333(.A1(G137gat), .A2(G154gat), .A3(G273gat), .A4(G290gat), .ZN(new_n462_));
  INV_X1    g0334(.A(new_n462_), .ZN(new_n463_));
  AOI22_X1  g0335(.A1(G137gat), .A2(G290gat), .B1(G154gat), .B2(G273gat), .ZN(new_n464_));
  OAI21_X1  g0336(.A(new_n379_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g0337(.A1(new_n382_), .A2(new_n462_), .ZN(new_n466_));
  NAND2_X1  g0338(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g0339(.A1(new_n300_), .A2(new_n150_), .ZN(new_n468_));
  OR2_X1    g0340(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g0341(.A1(new_n467_), .A2(new_n468_), .ZN(new_n470_));
  AOI21_X1  g0342(.A(new_n461_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g0343(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g0344(.A1(new_n469_), .A2(new_n470_), .A3(new_n461_), .ZN(new_n473_));
  AOI21_X1  g0345(.A(new_n460_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g0346(.A(new_n473_), .ZN(new_n475_));
  NOR3_X1   g0347(.A1(new_n475_), .A2(new_n471_), .A3(new_n459_), .ZN(new_n476_));
  OAI21_X1  g0348(.A(new_n458_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g0349(.A(new_n399_), .ZN(new_n478_));
  OAI21_X1  g0350(.A(new_n396_), .B1(new_n397_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g0351(.A1(new_n472_), .A2(new_n460_), .A3(new_n473_), .ZN(new_n480_));
  OAI21_X1  g0352(.A(new_n459_), .B1(new_n475_), .B2(new_n471_), .ZN(new_n481_));
  NAND3_X1  g0353(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NOR2_X1   g0354(.A1(new_n242_), .A2(new_n198_), .ZN(new_n483_));
  INV_X1    g0355(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g0356(.A1(new_n477_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g0357(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g0358(.A(new_n484_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n487_));
  NOR2_X1   g0359(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g0360(.A(new_n405_), .B1(new_n404_), .B2(new_n400_), .ZN(new_n489_));
  OAI21_X1  g0361(.A(new_n406_), .B1(new_n489_), .B2(new_n408_), .ZN(new_n490_));
  NAND2_X1  g0362(.A1(new_n490_), .A2(KEYINPUT12), .ZN(new_n491_));
  INV_X1    g0363(.A(KEYINPUT12), .ZN(new_n492_));
  OAI211_X1 g0364(.A(new_n492_), .B(new_n406_), .C1(new_n489_), .C2(new_n408_), .ZN(new_n493_));
  AOI21_X1  g0365(.A(new_n488_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g0366(.A(new_n492_), .B1(new_n411_), .B2(new_n406_), .ZN(new_n495_));
  INV_X1    g0367(.A(new_n487_), .ZN(new_n496_));
  NAND2_X1  g0368(.A1(new_n496_), .A2(new_n485_), .ZN(new_n497_));
  NOR2_X1   g0369(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g0370(.A1(new_n166_), .A2(new_n276_), .ZN(new_n499_));
  INV_X1    g0371(.A(new_n499_), .ZN(new_n500_));
  NOR3_X1   g0372(.A1(new_n494_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g0373(.A(new_n493_), .ZN(new_n502_));
  OAI21_X1  g0374(.A(new_n497_), .B1(new_n495_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g0375(.A1(new_n491_), .A2(new_n488_), .ZN(new_n504_));
  AOI21_X1  g0376(.A(new_n499_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g0377(.A(new_n457_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g0378(.A(new_n500_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n507_));
  NAND3_X1  g0379(.A1(new_n503_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n508_));
  OAI211_X1 g0380(.A(new_n507_), .B(new_n508_), .C1(new_n419_), .C2(new_n456_), .ZN(new_n509_));
  AOI21_X1  g0381(.A(new_n455_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g0382(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g0383(.A1(new_n506_), .A2(new_n509_), .A3(new_n455_), .ZN(new_n512_));
  AOI21_X1  g0384(.A(new_n453_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g0385(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g0386(.A1(new_n511_), .A2(new_n453_), .A3(new_n512_), .ZN(new_n515_));
  AOI21_X1  g0387(.A(new_n452_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g0388(.A(new_n515_), .ZN(new_n517_));
  NOR3_X1   g0389(.A1(new_n517_), .A2(new_n513_), .A3(new_n451_), .ZN(new_n518_));
  NOR2_X1   g0390(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g0391(.A1(new_n450_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g0392(.A(new_n434_), .B(new_n449_), .C1(new_n516_), .C2(new_n518_), .ZN(new_n521_));
  NAND2_X1  g0393(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g0394(.A1(new_n522_), .A2(G18gat), .A3(G409gat), .ZN(new_n523_));
  NAND2_X1  g0395(.A1(G18gat), .A2(G409gat), .ZN(new_n524_));
  NAND3_X1  g0396(.A1(new_n520_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n525_));
  NAND2_X1  g0397(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g0398(.A1(new_n448_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g0399(.A(new_n526_), .ZN(new_n528_));
  NOR3_X1   g0400(.A1(new_n440_), .A2(new_n439_), .A3(new_n368_), .ZN(new_n529_));
  OAI21_X1  g0401(.A(new_n441_), .B1(new_n529_), .B2(new_n444_), .ZN(new_n530_));
  NAND2_X1  g0402(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g0403(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g0404(.A(G426gat), .ZN(new_n533_));
  NOR2_X1   g0405(.A1(new_n129_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g0406(.A(new_n532_), .B(new_n534_), .ZN(G4241gat));
  NOR2_X1   g0407(.A1(new_n528_), .A2(new_n530_), .ZN(new_n536_));
  OAI21_X1  g0408(.A(new_n515_), .B1(new_n513_), .B2(new_n451_), .ZN(new_n537_));
  AND2_X1   g0409(.A1(new_n485_), .A2(new_n482_), .ZN(new_n538_));
  OAI21_X1  g0410(.A(new_n473_), .B1(new_n471_), .B2(new_n459_), .ZN(new_n539_));
  INV_X1    g0411(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g0412(.A1(new_n377_), .A2(new_n150_), .ZN(new_n541_));
  INV_X1    g0413(.A(G154gat), .ZN(new_n542_));
  INV_X1    g0414(.A(G171gat), .ZN(new_n543_));
  OAI22_X1  g0415(.A1(new_n542_), .A2(new_n133_), .B1(new_n543_), .B2(new_n130_), .ZN(new_n544_));
  NAND4_X1  g0416(.A1(G154gat), .A2(G171gat), .A3(G273gat), .A4(G290gat), .ZN(new_n545_));
  NAND3_X1  g0417(.A1(new_n544_), .A2(KEYINPUT13), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g0418(.A(KEYINPUT13), .ZN(new_n547_));
  OAI221_X1 g0419(.A(new_n547_), .B1(new_n542_), .B2(new_n133_), .C1(new_n543_), .C2(new_n130_), .ZN(new_n548_));
  NAND3_X1  g0420(.A1(new_n546_), .A2(new_n462_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g0421(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g0422(.A(new_n462_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n551_));
  OAI21_X1  g0423(.A(new_n541_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g0424(.A1(new_n465_), .A2(new_n468_), .ZN(new_n553_));
  NAND2_X1  g0425(.A1(new_n553_), .A2(new_n466_), .ZN(new_n554_));
  INV_X1    g0426(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g0427(.A1(new_n546_), .A2(new_n548_), .ZN(new_n556_));
  NAND2_X1  g0428(.A1(new_n556_), .A2(new_n463_), .ZN(new_n557_));
  INV_X1    g0429(.A(new_n541_), .ZN(new_n558_));
  NAND3_X1  g0430(.A1(new_n557_), .A2(new_n558_), .A3(new_n549_), .ZN(new_n559_));
  NAND3_X1  g0431(.A1(new_n552_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g0432(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g0433(.A(new_n555_), .B1(new_n552_), .B2(new_n559_), .ZN(new_n562_));
  NOR2_X1   g0434(.A1(new_n300_), .A2(new_n159_), .ZN(new_n563_));
  NOR3_X1   g0435(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g0436(.A(new_n563_), .ZN(new_n565_));
  NOR3_X1   g0437(.A1(new_n550_), .A2(new_n551_), .A3(new_n541_), .ZN(new_n566_));
  AOI21_X1  g0438(.A(new_n558_), .B1(new_n557_), .B2(new_n549_), .ZN(new_n567_));
  OAI21_X1  g0439(.A(new_n554_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g0440(.A(new_n565_), .B1(new_n568_), .B2(new_n560_), .ZN(new_n569_));
  OAI21_X1  g0441(.A(new_n540_), .B1(new_n564_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g0442(.A1(new_n243_), .A2(new_n198_), .ZN(new_n571_));
  INV_X1    g0443(.A(new_n571_), .ZN(new_n572_));
  OAI21_X1  g0444(.A(new_n563_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n573_));
  NAND3_X1  g0445(.A1(new_n568_), .A2(new_n565_), .A3(new_n560_), .ZN(new_n574_));
  NAND3_X1  g0446(.A1(new_n573_), .A2(new_n539_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g0447(.A1(new_n570_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g0448(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g0449(.A(new_n572_), .B1(new_n570_), .B2(new_n575_), .ZN(new_n578_));
  OAI21_X1  g0450(.A(new_n538_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g0451(.A1(new_n485_), .A2(new_n482_), .ZN(new_n580_));
  NOR3_X1   g0452(.A1(new_n564_), .A2(new_n569_), .A3(new_n540_), .ZN(new_n581_));
  AOI21_X1  g0453(.A(new_n539_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n582_));
  OAI21_X1  g0454(.A(new_n571_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g0455(.A1(new_n580_), .A2(new_n583_), .A3(new_n576_), .ZN(new_n584_));
  NAND2_X1  g0456(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g0457(.A1(new_n242_), .A2(new_n276_), .ZN(new_n586_));
  INV_X1    g0458(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g0459(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g0460(.A1(new_n579_), .A2(new_n586_), .A3(new_n584_), .ZN(new_n589_));
  AND2_X1   g0461(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g0462(.A1(new_n488_), .A2(new_n490_), .ZN(new_n591_));
  INV_X1    g0463(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g0464(.A1(new_n505_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g0465(.A(KEYINPUT14), .ZN(new_n594_));
  AOI21_X1  g0466(.A(new_n594_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n595_));
  OAI21_X1  g0467(.A(new_n590_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g0468(.A1(new_n166_), .A2(new_n289_), .ZN(new_n597_));
  INV_X1    g0469(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g0470(.A1(new_n507_), .A2(new_n591_), .ZN(new_n599_));
  INV_X1    g0471(.A(new_n595_), .ZN(new_n600_));
  NAND2_X1  g0472(.A1(new_n588_), .A2(new_n589_), .ZN(new_n601_));
  NAND3_X1  g0473(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g0474(.A1(new_n596_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g0475(.A(new_n602_), .ZN(new_n604_));
  AOI21_X1  g0476(.A(new_n601_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n605_));
  OAI21_X1  g0477(.A(new_n597_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g0478(.A(KEYINPUT15), .ZN(new_n607_));
  AND3_X1   g0479(.A1(new_n512_), .A2(new_n607_), .A3(new_n509_), .ZN(new_n608_));
  AOI21_X1  g0480(.A(new_n607_), .B1(new_n512_), .B2(new_n509_), .ZN(new_n609_));
  OAI211_X1 g0481(.A(new_n603_), .B(new_n606_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g0482(.A1(new_n457_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n611_));
  AOI21_X1  g0483(.A(new_n611_), .B1(new_n455_), .B2(new_n506_), .ZN(new_n612_));
  NAND2_X1  g0484(.A1(new_n612_), .A2(new_n607_), .ZN(new_n613_));
  INV_X1    g0485(.A(new_n603_), .ZN(new_n614_));
  AOI21_X1  g0486(.A(new_n598_), .B1(new_n596_), .B2(new_n602_), .ZN(new_n615_));
  OAI21_X1  g0487(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g0488(.A1(new_n610_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g0489(.A1(new_n165_), .A2(new_n363_), .ZN(new_n618_));
  INV_X1    g0490(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g0491(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g0492(.A1(new_n610_), .A2(new_n618_), .A3(new_n616_), .ZN(new_n621_));
  AOI21_X1  g0493(.A(new_n537_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g0494(.A(new_n622_), .ZN(new_n623_));
  NAND3_X1  g0495(.A1(new_n620_), .A2(new_n537_), .A3(new_n621_), .ZN(new_n624_));
  NOR2_X1   g0496(.A1(new_n218_), .A2(new_n443_), .ZN(new_n625_));
  INV_X1    g0497(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g0498(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g0499(.A(new_n621_), .ZN(new_n628_));
  INV_X1    g0500(.A(new_n537_), .ZN(new_n629_));
  AOI21_X1  g0501(.A(new_n618_), .B1(new_n610_), .B2(new_n616_), .ZN(new_n630_));
  NOR3_X1   g0502(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g0503(.A(new_n625_), .B1(new_n631_), .B2(new_n622_), .ZN(new_n632_));
  NAND2_X1  g0504(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g0505(.A1(new_n633_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n634_));
  NAND2_X1  g0506(.A1(new_n525_), .A2(new_n520_), .ZN(new_n635_));
  NAND3_X1  g0507(.A1(new_n635_), .A2(new_n627_), .A3(new_n632_), .ZN(new_n636_));
  NOR2_X1   g0508(.A1(new_n132_), .A2(new_n533_), .ZN(new_n637_));
  INV_X1    g0509(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g0510(.A1(new_n634_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g0511(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g0512(.A(new_n638_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n641_));
  OAI221_X1 g0513(.A(new_n531_), .B1(new_n536_), .B2(new_n534_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g0514(.A(new_n531_), .B1(new_n536_), .B2(new_n534_), .ZN(new_n643_));
  INV_X1    g0515(.A(new_n641_), .ZN(new_n644_));
  NAND3_X1  g0516(.A1(new_n643_), .A2(new_n644_), .A3(new_n639_), .ZN(new_n645_));
  AND3_X1   g0517(.A1(new_n642_), .A2(new_n645_), .A3(KEYINPUT16), .ZN(new_n646_));
  AOI21_X1  g0518(.A(KEYINPUT16), .B1(new_n642_), .B2(new_n645_), .ZN(new_n647_));
  INV_X1    g0519(.A(G443gat), .ZN(new_n648_));
  NOR2_X1   g0520(.A1(new_n129_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g0521(.A(new_n649_), .ZN(new_n650_));
  OR3_X1    g0522(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g0523(.A(new_n650_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n652_));
  NAND2_X1  g0524(.A1(new_n651_), .A2(new_n652_), .ZN(G4591gat));
  INV_X1    g0525(.A(G460gat), .ZN(new_n654_));
  NOR2_X1   g0526(.A1(new_n129_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g0527(.A1(new_n639_), .A2(new_n636_), .ZN(new_n656_));
  NOR2_X1   g0528(.A1(new_n218_), .A2(new_n533_), .ZN(new_n657_));
  NOR3_X1   g0529(.A1(new_n614_), .A2(new_n615_), .A3(new_n612_), .ZN(new_n658_));
  NOR2_X1   g0530(.A1(new_n630_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g0531(.A1(new_n599_), .A2(new_n601_), .ZN(new_n660_));
  NAND2_X1  g0532(.A1(new_n603_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0533(.A1(new_n584_), .A2(new_n586_), .ZN(new_n662_));
  NAND2_X1  g0534(.A1(new_n662_), .A2(new_n579_), .ZN(new_n663_));
  INV_X1    g0535(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g0536(.A1(new_n243_), .A2(new_n276_), .ZN(new_n665_));
  INV_X1    g0537(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g0538(.A1(G154gat), .A2(G307gat), .ZN(new_n667_));
  INV_X1    g0539(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g0540(.A1(G188gat), .A2(G273gat), .ZN(new_n669_));
  OAI21_X1  g0541(.A(new_n669_), .B1(new_n543_), .B2(new_n133_), .ZN(new_n670_));
  NAND4_X1  g0542(.A1(G171gat), .A2(G188gat), .A3(G273gat), .A4(G290gat), .ZN(new_n671_));
  NOR2_X1   g0543(.A1(new_n542_), .A2(new_n133_), .ZN(new_n672_));
  NOR2_X1   g0544(.A1(new_n543_), .A2(new_n130_), .ZN(new_n673_));
  AOI22_X1  g0545(.A1(new_n670_), .A2(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g0546(.A(new_n671_), .ZN(new_n675_));
  NOR2_X1   g0547(.A1(new_n675_), .A2(new_n545_), .ZN(new_n676_));
  OAI21_X1  g0548(.A(new_n668_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g0549(.A1(new_n670_), .A2(new_n671_), .ZN(new_n678_));
  NAND2_X1  g0550(.A1(new_n678_), .A2(new_n545_), .ZN(new_n679_));
  NAND3_X1  g0551(.A1(new_n672_), .A2(new_n673_), .A3(new_n671_), .ZN(new_n680_));
  NAND3_X1  g0552(.A1(new_n679_), .A2(new_n667_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g0553(.A1(new_n677_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g0554(.A1(new_n559_), .A2(new_n682_), .A3(new_n549_), .ZN(new_n683_));
  NOR2_X1   g0555(.A1(new_n377_), .A2(new_n159_), .ZN(new_n684_));
  INV_X1    g0556(.A(new_n684_), .ZN(new_n685_));
  AND2_X1   g0557(.A1(new_n677_), .A2(new_n681_), .ZN(new_n686_));
  OAI21_X1  g0558(.A(new_n549_), .B1(new_n551_), .B2(new_n541_), .ZN(new_n687_));
  NAND2_X1  g0559(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND3_X1   g0560(.A1(new_n683_), .A2(new_n685_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g0561(.A(new_n685_), .B1(new_n683_), .B2(new_n688_), .ZN(new_n690_));
  OAI211_X1 g0562(.A(new_n574_), .B(new_n560_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g0563(.A1(new_n683_), .A2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g0564(.A1(new_n692_), .A2(new_n684_), .ZN(new_n693_));
  OAI21_X1  g0565(.A(new_n560_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n694_));
  NAND3_X1  g0566(.A1(new_n683_), .A2(new_n688_), .A3(new_n685_), .ZN(new_n695_));
  NAND3_X1  g0567(.A1(new_n693_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g0568(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g0569(.A1(new_n300_), .A2(new_n198_), .ZN(new_n698_));
  INV_X1    g0570(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g0571(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g0572(.A(KEYINPUT17), .ZN(new_n701_));
  NAND2_X1  g0573(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g0574(.A1(new_n691_), .A2(new_n698_), .A3(new_n696_), .ZN(new_n703_));
  NAND2_X1  g0575(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g0576(.A1(new_n576_), .A2(new_n575_), .ZN(new_n705_));
  NAND3_X1  g0577(.A1(new_n702_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g0578(.A(new_n581_), .B1(new_n572_), .B2(new_n570_), .ZN(new_n707_));
  OAI211_X1 g0579(.A(new_n700_), .B(new_n703_), .C1(new_n707_), .C2(new_n701_), .ZN(new_n708_));
  AOI21_X1  g0580(.A(new_n666_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g0581(.A(new_n709_), .ZN(new_n710_));
  NAND3_X1  g0582(.A1(new_n706_), .A2(new_n708_), .A3(new_n666_), .ZN(new_n711_));
  AOI21_X1  g0583(.A(new_n664_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g0584(.A(new_n711_), .ZN(new_n713_));
  NOR3_X1   g0585(.A1(new_n713_), .A2(new_n709_), .A3(new_n663_), .ZN(new_n714_));
  NOR2_X1   g0586(.A1(new_n242_), .A2(new_n289_), .ZN(new_n715_));
  NOR3_X1   g0587(.A1(new_n712_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g0588(.A(new_n715_), .ZN(new_n717_));
  OAI21_X1  g0589(.A(new_n663_), .B1(new_n713_), .B2(new_n709_), .ZN(new_n718_));
  NAND3_X1  g0590(.A1(new_n710_), .A2(new_n664_), .A3(new_n711_), .ZN(new_n719_));
  AOI21_X1  g0591(.A(new_n717_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g0592(.A1(new_n716_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g0593(.A1(new_n661_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g0594(.A(new_n603_), .B(new_n660_), .C1(new_n716_), .C2(new_n720_), .ZN(new_n723_));
  NAND2_X1  g0595(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g0596(.A1(new_n166_), .A2(new_n363_), .ZN(new_n725_));
  NAND2_X1  g0597(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g0598(.A(new_n725_), .ZN(new_n727_));
  NAND3_X1  g0599(.A1(new_n722_), .A2(new_n727_), .A3(new_n723_), .ZN(new_n728_));
  NAND2_X1  g0600(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g0601(.A1(new_n659_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g0602(.A(new_n728_), .B(new_n726_), .C1(new_n630_), .C2(new_n658_), .ZN(new_n731_));
  NAND2_X1  g0603(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g0604(.A1(new_n165_), .A2(new_n443_), .ZN(new_n733_));
  NAND2_X1  g0605(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g0606(.A(new_n624_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n735_));
  INV_X1    g0607(.A(new_n733_), .ZN(new_n736_));
  NAND3_X1  g0608(.A1(new_n730_), .A2(new_n736_), .A3(new_n731_), .ZN(new_n737_));
  NAND3_X1  g0609(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g0610(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g0611(.A(new_n735_), .B1(new_n734_), .B2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g0612(.A(new_n657_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g0613(.A(new_n735_), .ZN(new_n742_));
  INV_X1    g0614(.A(new_n737_), .ZN(new_n743_));
  AOI21_X1  g0615(.A(new_n736_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n744_));
  OAI21_X1  g0616(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g0617(.A(new_n657_), .ZN(new_n746_));
  NAND3_X1  g0618(.A1(new_n745_), .A2(new_n746_), .A3(new_n738_), .ZN(new_n747_));
  AOI21_X1  g0619(.A(new_n656_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g0620(.A(new_n748_), .ZN(new_n749_));
  NAND3_X1  g0621(.A1(new_n656_), .A2(new_n747_), .A3(new_n741_), .ZN(new_n750_));
  NAND2_X1  g0622(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g0623(.A1(new_n132_), .A2(new_n648_), .ZN(new_n752_));
  INV_X1    g0624(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g0625(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g0626(.A1(new_n749_), .A2(new_n752_), .A3(new_n750_), .ZN(new_n755_));
  NAND2_X1  g0627(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g0628(.A1(new_n756_), .A2(new_n652_), .A3(new_n645_), .ZN(new_n757_));
  NAND2_X1  g0629(.A1(new_n755_), .A2(KEYINPUT18), .ZN(new_n758_));
  NAND2_X1  g0630(.A1(new_n645_), .A2(new_n649_), .ZN(new_n759_));
  AND2_X1   g0631(.A1(new_n759_), .A2(new_n642_), .ZN(new_n760_));
  INV_X1    g0632(.A(KEYINPUT18), .ZN(new_n761_));
  NAND4_X1  g0633(.A1(new_n749_), .A2(new_n761_), .A3(new_n752_), .A4(new_n750_), .ZN(new_n762_));
  NAND4_X1  g0634(.A1(new_n758_), .A2(new_n760_), .A3(new_n754_), .A4(new_n762_), .ZN(new_n763_));
  AOI21_X1  g0635(.A(new_n655_), .B1(new_n757_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g0636(.A(new_n764_), .ZN(new_n765_));
  NAND3_X1  g0637(.A1(new_n757_), .A2(new_n655_), .A3(new_n763_), .ZN(new_n766_));
  NAND2_X1  g0638(.A1(new_n765_), .A2(new_n766_), .ZN(G4946gat));
  NAND2_X1  g0639(.A1(new_n750_), .A2(new_n752_), .ZN(new_n768_));
  NAND2_X1  g0640(.A1(new_n749_), .A2(new_n768_), .ZN(new_n769_));
  AND2_X1   g0641(.A1(new_n659_), .A2(new_n729_), .ZN(new_n770_));
  OAI21_X1  g0642(.A(new_n731_), .B1(new_n770_), .B2(new_n733_), .ZN(new_n771_));
  INV_X1    g0643(.A(new_n723_), .ZN(new_n772_));
  OAI21_X1  g0644(.A(new_n722_), .B1(new_n772_), .B2(new_n725_), .ZN(new_n773_));
  NAND2_X1  g0645(.A1(G86gat), .A2(G392gat), .ZN(new_n774_));
  XNOR2_X1  g0646(.A(new_n774_), .B(KEYINPUT21), .ZN(new_n775_));
  INV_X1    g0647(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g0648(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n777_));
  NAND2_X1  g0649(.A1(new_n704_), .A2(new_n705_), .ZN(new_n778_));
  NAND2_X1  g0650(.A1(new_n711_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g0651(.A1(new_n300_), .A2(new_n276_), .ZN(new_n780_));
  NAND2_X1  g0652(.A1(new_n696_), .A2(new_n698_), .ZN(new_n781_));
  NAND2_X1  g0653(.A1(new_n781_), .A2(new_n691_), .ZN(new_n782_));
  NAND2_X1  g0654(.A1(G188gat), .A2(G290gat), .ZN(new_n783_));
  NAND2_X1  g0655(.A1(G205gat), .A2(G273gat), .ZN(new_n784_));
  NAND2_X1  g0656(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g0657(.A1(G188gat), .A2(G205gat), .A3(G273gat), .A4(G290gat), .ZN(new_n786_));
  NAND2_X1  g0658(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g0659(.A1(new_n787_), .A2(new_n671_), .ZN(new_n788_));
  NAND2_X1  g0660(.A1(new_n675_), .A2(new_n786_), .ZN(new_n789_));
  NAND2_X1  g0661(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g0662(.A1(G171gat), .A2(G307gat), .ZN(new_n791_));
  INV_X1    g0663(.A(KEYINPUT19), .ZN(new_n792_));
  NAND2_X1  g0664(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g0665(.A1(KEYINPUT19), .A2(G171gat), .A3(G307gat), .ZN(new_n794_));
  NAND2_X1  g0666(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g0667(.A(KEYINPUT20), .ZN(new_n796_));
  NAND2_X1  g0668(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g0669(.A1(new_n793_), .A2(KEYINPUT20), .A3(new_n794_), .ZN(new_n798_));
  NAND2_X1  g0670(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g0671(.A1(new_n790_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g0672(.A(new_n674_), .B1(new_n667_), .B2(new_n680_), .ZN(new_n801_));
  NAND3_X1  g0673(.A1(new_n788_), .A2(new_n789_), .A3(new_n798_), .ZN(new_n802_));
  NAND3_X1  g0674(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g0675(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g0676(.A(new_n801_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n805_));
  NOR2_X1   g0677(.A1(new_n542_), .A2(new_n159_), .ZN(new_n806_));
  NOR3_X1   g0678(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g0679(.A(new_n806_), .ZN(new_n808_));
  NAND2_X1  g0680(.A1(new_n800_), .A2(new_n802_), .ZN(new_n809_));
  INV_X1    g0681(.A(new_n801_), .ZN(new_n810_));
  NAND2_X1  g0682(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g0683(.A(new_n808_), .B1(new_n811_), .B2(new_n803_), .ZN(new_n812_));
  OAI211_X1 g0684(.A(new_n688_), .B(new_n695_), .C1(new_n807_), .C2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g0685(.A1(new_n377_), .A2(new_n198_), .ZN(new_n814_));
  INV_X1    g0686(.A(new_n814_), .ZN(new_n815_));
  NOR2_X1   g0687(.A1(new_n686_), .A2(new_n687_), .ZN(new_n816_));
  OAI21_X1  g0688(.A(new_n688_), .B1(new_n816_), .B2(new_n684_), .ZN(new_n817_));
  OAI21_X1  g0689(.A(new_n806_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n818_));
  NAND3_X1  g0690(.A1(new_n811_), .A2(new_n808_), .A3(new_n803_), .ZN(new_n819_));
  NAND3_X1  g0691(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  AND3_X1   g0692(.A1(new_n813_), .A2(new_n815_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g0693(.A(new_n815_), .B1(new_n813_), .B2(new_n820_), .ZN(new_n822_));
  NOR3_X1   g0694(.A1(new_n782_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g0695(.A1(new_n813_), .A2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g0696(.A1(new_n824_), .A2(new_n814_), .ZN(new_n825_));
  NAND3_X1  g0697(.A1(new_n813_), .A2(new_n815_), .A3(new_n820_), .ZN(new_n826_));
  AOI22_X1  g0698(.A1(new_n825_), .A2(new_n826_), .B1(new_n691_), .B2(new_n781_), .ZN(new_n827_));
  OAI21_X1  g0699(.A(new_n780_), .B1(new_n823_), .B2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g0700(.A1(new_n825_), .A2(new_n691_), .A3(new_n826_), .A4(new_n781_), .ZN(new_n829_));
  NOR2_X1   g0701(.A1(new_n689_), .A2(new_n690_), .ZN(new_n830_));
  AOI21_X1  g0702(.A(new_n699_), .B1(new_n830_), .B2(new_n694_), .ZN(new_n831_));
  AOI21_X1  g0703(.A(new_n694_), .B1(new_n695_), .B2(new_n693_), .ZN(new_n832_));
  OAI22_X1  g0704(.A1(new_n821_), .A2(new_n822_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g0705(.A(new_n780_), .ZN(new_n834_));
  NAND3_X1  g0706(.A1(new_n829_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AND2_X1   g0707(.A1(new_n828_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g0708(.A1(new_n779_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g0709(.A1(new_n243_), .A2(new_n289_), .ZN(new_n838_));
  INV_X1    g0710(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g0711(.A1(new_n828_), .A2(new_n835_), .ZN(new_n840_));
  NAND3_X1  g0712(.A1(new_n840_), .A2(new_n711_), .A3(new_n778_), .ZN(new_n841_));
  NAND3_X1  g0713(.A1(new_n837_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g0714(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g0715(.A(new_n839_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n844_));
  OAI21_X1  g0716(.A(new_n777_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g0717(.A(new_n844_), .ZN(new_n846_));
  OAI21_X1  g0718(.A(new_n719_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n847_));
  NAND3_X1  g0719(.A1(new_n846_), .A2(new_n847_), .A3(new_n842_), .ZN(new_n848_));
  AOI21_X1  g0720(.A(new_n776_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g0721(.A(new_n849_), .ZN(new_n850_));
  NAND3_X1  g0722(.A1(new_n845_), .A2(new_n848_), .A3(new_n774_), .ZN(new_n851_));
  NAND3_X1  g0723(.A1(new_n773_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AND3_X1   g0724(.A1(new_n845_), .A2(new_n848_), .A3(new_n776_), .ZN(new_n853_));
  OAI211_X1 g0725(.A(new_n728_), .B(new_n722_), .C1(new_n853_), .C2(new_n849_), .ZN(new_n854_));
  NAND2_X1  g0726(.A1(G69gat), .A2(G409gat), .ZN(new_n855_));
  AND3_X1   g0727(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g0728(.A(new_n855_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n857_));
  NOR2_X1   g0729(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g0730(.A1(new_n771_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g0731(.A(new_n737_), .B(new_n731_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n860_));
  NOR2_X1   g0732(.A1(new_n165_), .A2(new_n533_), .ZN(new_n861_));
  INV_X1    g0733(.A(new_n861_), .ZN(new_n862_));
  AND3_X1   g0734(.A1(new_n859_), .A2(new_n860_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g0735(.A(new_n862_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n864_));
  OAI211_X1 g0736(.A(new_n747_), .B(new_n738_), .C1(new_n863_), .C2(new_n864_), .ZN(new_n865_));
  AND2_X1   g0737(.A1(new_n771_), .A2(new_n858_), .ZN(new_n866_));
  NOR2_X1   g0738(.A1(new_n771_), .A2(new_n858_), .ZN(new_n867_));
  OAI21_X1  g0739(.A(new_n861_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g0740(.A(new_n738_), .B1(new_n740_), .B2(new_n657_), .ZN(new_n869_));
  NAND3_X1  g0741(.A1(new_n859_), .A2(new_n860_), .A3(new_n862_), .ZN(new_n870_));
  NAND3_X1  g0742(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  NAND2_X1  g0743(.A1(G35gat), .A2(G443gat), .ZN(new_n872_));
  NAND3_X1  g0744(.A1(new_n865_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g0745(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g0746(.A(new_n872_), .B1(new_n865_), .B2(new_n871_), .ZN(new_n875_));
  OAI21_X1  g0747(.A(new_n769_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g0748(.A1(G18gat), .A2(G460gat), .ZN(new_n877_));
  INV_X1    g0749(.A(new_n875_), .ZN(new_n878_));
  NAND4_X1  g0750(.A1(new_n768_), .A2(new_n749_), .A3(new_n878_), .A4(new_n873_), .ZN(new_n879_));
  NAND3_X1  g0751(.A1(new_n876_), .A2(new_n877_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g0752(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g0753(.A(new_n877_), .B1(new_n876_), .B2(new_n879_), .ZN(new_n882_));
  NOR2_X1   g0754(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g0755(.A1(new_n756_), .A2(new_n760_), .ZN(new_n884_));
  INV_X1    g0756(.A(new_n884_), .ZN(new_n885_));
  NOR3_X1   g0757(.A1(new_n764_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g0758(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g0759(.A(new_n883_), .B1(new_n764_), .B2(new_n885_), .ZN(new_n888_));
  NAND2_X1  g0760(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g0761(.A(G477gat), .ZN(new_n890_));
  NOR2_X1   g0762(.A1(new_n129_), .A2(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g0763(.A(new_n889_), .B(new_n891_), .ZN(G5308gat));
  OAI21_X1  g0764(.A(new_n888_), .B1(new_n886_), .B2(new_n891_), .ZN(new_n893_));
  NAND2_X1  g0765(.A1(new_n880_), .A2(new_n879_), .ZN(new_n894_));
  NAND2_X1  g0766(.A1(new_n873_), .A2(KEYINPUT22), .ZN(new_n895_));
  NOR2_X1   g0767(.A1(new_n166_), .A2(new_n533_), .ZN(new_n896_));
  NOR2_X1   g0768(.A1(new_n300_), .A2(new_n289_), .ZN(new_n897_));
  NOR2_X1   g0769(.A1(new_n377_), .A2(new_n276_), .ZN(new_n898_));
  NOR2_X1   g0770(.A1(new_n542_), .A2(new_n198_), .ZN(new_n899_));
  XNOR2_X1  g0771(.A(new_n899_), .B(KEYINPUT28), .ZN(new_n900_));
  NAND2_X1  g0772(.A1(G205gat), .A2(G290gat), .ZN(new_n901_));
  NAND2_X1  g0773(.A1(G222gat), .A2(G273gat), .ZN(new_n902_));
  INV_X1    g0774(.A(KEYINPUT26), .ZN(new_n903_));
  AND3_X1   g0775(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g0776(.A(new_n901_), .B1(new_n903_), .B2(new_n902_), .ZN(new_n905_));
  OAI21_X1  g0777(.A(new_n786_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  NAND4_X1  g0778(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n907_));
  INV_X1    g0779(.A(new_n907_), .ZN(new_n908_));
  OR2_X1    g0780(.A1(new_n908_), .A2(new_n786_), .ZN(new_n909_));
  NAND2_X1  g0781(.A1(new_n906_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g0782(.A1(G188gat), .A2(G307gat), .ZN(new_n911_));
  INV_X1    g0783(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g0784(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  AND2_X1   g0785(.A1(new_n793_), .A2(new_n794_), .ZN(new_n914_));
  AOI22_X1  g0786(.A1(new_n914_), .A2(new_n789_), .B1(new_n787_), .B2(new_n671_), .ZN(new_n915_));
  NAND3_X1  g0787(.A1(new_n906_), .A2(new_n911_), .A3(new_n909_), .ZN(new_n916_));
  NAND3_X1  g0788(.A1(new_n913_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g0789(.A(KEYINPUT27), .ZN(new_n918_));
  NAND2_X1  g0790(.A1(new_n901_), .A2(new_n902_), .ZN(new_n919_));
  NAND3_X1  g0791(.A1(new_n919_), .A2(new_n786_), .A3(new_n907_), .ZN(new_n920_));
  INV_X1    g0792(.A(KEYINPUT25), .ZN(new_n921_));
  NAND2_X1  g0793(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND4_X1  g0794(.A1(new_n919_), .A2(KEYINPUT25), .A3(new_n786_), .A4(new_n907_), .ZN(new_n923_));
  NAND3_X1  g0795(.A1(new_n905_), .A2(G188gat), .A3(G273gat), .ZN(new_n924_));
  NAND4_X1  g0796(.A1(new_n922_), .A2(new_n912_), .A3(new_n923_), .A4(new_n924_), .ZN(new_n925_));
  NAND2_X1  g0797(.A1(new_n925_), .A2(new_n916_), .ZN(new_n926_));
  INV_X1    g0798(.A(new_n915_), .ZN(new_n927_));
  AOI21_X1  g0799(.A(new_n918_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  AOI211_X1 g0800(.A(KEYINPUT27), .B(new_n915_), .C1(new_n925_), .C2(new_n916_), .ZN(new_n929_));
  OAI21_X1  g0801(.A(new_n917_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g0802(.A1(new_n543_), .A2(new_n159_), .ZN(new_n931_));
  INV_X1    g0803(.A(new_n931_), .ZN(new_n932_));
  NAND2_X1  g0804(.A1(new_n930_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g0805(.A1(new_n819_), .A2(new_n811_), .ZN(new_n934_));
  OAI211_X1 g0806(.A(new_n931_), .B(new_n917_), .C1(new_n928_), .C2(new_n929_), .ZN(new_n935_));
  AND3_X1   g0807(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  AOI21_X1  g0808(.A(new_n934_), .B1(new_n933_), .B2(new_n935_), .ZN(new_n937_));
  OAI21_X1  g0809(.A(new_n900_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g0810(.A1(new_n826_), .A2(new_n820_), .ZN(new_n939_));
  INV_X1    g0811(.A(new_n934_), .ZN(new_n940_));
  NAND2_X1  g0812(.A1(new_n926_), .A2(new_n927_), .ZN(new_n941_));
  NAND2_X1  g0813(.A1(new_n941_), .A2(KEYINPUT27), .ZN(new_n942_));
  NAND3_X1  g0814(.A1(new_n926_), .A2(new_n918_), .A3(new_n927_), .ZN(new_n943_));
  NAND2_X1  g0815(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g0816(.A(new_n931_), .B1(new_n944_), .B2(new_n917_), .ZN(new_n945_));
  INV_X1    g0817(.A(new_n935_), .ZN(new_n946_));
  OAI21_X1  g0818(.A(new_n940_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  NAND3_X1  g0819(.A1(new_n933_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n948_));
  INV_X1    g0820(.A(new_n899_), .ZN(new_n949_));
  NAND3_X1  g0821(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AND3_X1   g0822(.A1(new_n938_), .A2(new_n939_), .A3(new_n950_), .ZN(new_n951_));
  INV_X1    g0823(.A(new_n900_), .ZN(new_n952_));
  NAND3_X1  g0824(.A1(new_n947_), .A2(new_n948_), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g0825(.A(new_n939_), .B1(new_n938_), .B2(new_n953_), .ZN(new_n954_));
  OAI21_X1  g0826(.A(new_n898_), .B1(new_n951_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g0827(.A(new_n939_), .ZN(new_n956_));
  NOR3_X1   g0828(.A1(new_n936_), .A2(new_n937_), .A3(new_n900_), .ZN(new_n957_));
  AOI21_X1  g0829(.A(new_n952_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n958_));
  OAI21_X1  g0830(.A(new_n956_), .B1(new_n957_), .B2(new_n958_), .ZN(new_n959_));
  INV_X1    g0831(.A(new_n898_), .ZN(new_n960_));
  NAND3_X1  g0832(.A1(new_n938_), .A2(new_n939_), .A3(new_n950_), .ZN(new_n961_));
  NAND3_X1  g0833(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(new_n962_));
  INV_X1    g0834(.A(KEYINPUT24), .ZN(new_n963_));
  OAI21_X1  g0835(.A(new_n963_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n964_));
  NAND3_X1  g0836(.A1(new_n825_), .A2(KEYINPUT24), .A3(new_n826_), .ZN(new_n965_));
  INV_X1    g0837(.A(new_n782_), .ZN(new_n966_));
  NAND3_X1  g0838(.A1(new_n964_), .A2(new_n965_), .A3(new_n966_), .ZN(new_n967_));
  NAND2_X1  g0839(.A1(new_n835_), .A2(new_n967_), .ZN(new_n968_));
  AND3_X1   g0840(.A1(new_n955_), .A2(new_n962_), .A3(new_n968_), .ZN(new_n969_));
  AOI21_X1  g0841(.A(new_n968_), .B1(new_n955_), .B2(new_n962_), .ZN(new_n970_));
  OAI21_X1  g0842(.A(new_n897_), .B1(new_n969_), .B2(new_n970_), .ZN(new_n971_));
  INV_X1    g0843(.A(KEYINPUT23), .ZN(new_n972_));
  NAND2_X1  g0844(.A1(new_n837_), .A2(new_n972_), .ZN(new_n973_));
  AND2_X1   g0845(.A1(new_n835_), .A2(new_n967_), .ZN(new_n974_));
  NOR3_X1   g0846(.A1(new_n951_), .A2(new_n954_), .A3(new_n898_), .ZN(new_n975_));
  AOI21_X1  g0847(.A(new_n960_), .B1(new_n959_), .B2(new_n961_), .ZN(new_n976_));
  OAI21_X1  g0848(.A(new_n974_), .B1(new_n975_), .B2(new_n976_), .ZN(new_n977_));
  INV_X1    g0849(.A(new_n897_), .ZN(new_n978_));
  NAND3_X1  g0850(.A1(new_n955_), .A2(new_n968_), .A3(new_n962_), .ZN(new_n979_));
  NAND3_X1  g0851(.A1(new_n977_), .A2(new_n978_), .A3(new_n979_), .ZN(new_n980_));
  NAND3_X1  g0852(.A1(new_n971_), .A2(new_n973_), .A3(new_n980_), .ZN(new_n981_));
  AOI21_X1  g0853(.A(new_n840_), .B1(new_n711_), .B2(new_n778_), .ZN(new_n982_));
  AOI21_X1  g0854(.A(new_n982_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n983_));
  NAND2_X1  g0855(.A1(new_n981_), .A2(new_n983_), .ZN(new_n984_));
  INV_X1    g0856(.A(new_n841_), .ZN(new_n985_));
  OAI21_X1  g0857(.A(new_n837_), .B1(new_n985_), .B2(new_n838_), .ZN(new_n986_));
  NAND4_X1  g0858(.A1(new_n986_), .A2(new_n973_), .A3(new_n971_), .A4(new_n980_), .ZN(new_n987_));
  NAND2_X1  g0859(.A1(new_n984_), .A2(new_n987_), .ZN(new_n988_));
  INV_X1    g0860(.A(KEYINPUT29), .ZN(new_n989_));
  NAND2_X1  g0861(.A1(new_n988_), .A2(new_n989_), .ZN(new_n990_));
  NAND2_X1  g0862(.A1(G103gat), .A2(G392gat), .ZN(new_n991_));
  NAND3_X1  g0863(.A1(new_n984_), .A2(new_n987_), .A3(KEYINPUT29), .ZN(new_n992_));
  NAND3_X1  g0864(.A1(new_n990_), .A2(new_n991_), .A3(new_n992_), .ZN(new_n993_));
  INV_X1    g0865(.A(new_n848_), .ZN(new_n994_));
  AOI21_X1  g0866(.A(new_n994_), .B1(new_n845_), .B2(new_n776_), .ZN(new_n995_));
  NAND4_X1  g0867(.A1(new_n988_), .A2(new_n989_), .A3(G103gat), .A4(G392gat), .ZN(new_n996_));
  NAND3_X1  g0868(.A1(new_n993_), .A2(new_n995_), .A3(new_n996_), .ZN(new_n997_));
  INV_X1    g0869(.A(KEYINPUT30), .ZN(new_n998_));
  NAND2_X1  g0870(.A1(new_n997_), .A2(new_n998_), .ZN(new_n999_));
  NAND4_X1  g0871(.A1(new_n993_), .A2(KEYINPUT30), .A3(new_n995_), .A4(new_n996_), .ZN(new_n1000_));
  NAND2_X1  g0872(.A1(new_n993_), .A2(new_n996_), .ZN(new_n1001_));
  NAND2_X1  g0873(.A1(new_n851_), .A2(new_n848_), .ZN(new_n1002_));
  NAND2_X1  g0874(.A1(new_n1001_), .A2(new_n1002_), .ZN(new_n1003_));
  NAND3_X1  g0875(.A1(new_n999_), .A2(new_n1000_), .A3(new_n1003_), .ZN(new_n1004_));
  NOR2_X1   g0876(.A1(new_n242_), .A2(new_n443_), .ZN(new_n1005_));
  INV_X1    g0877(.A(new_n1005_), .ZN(new_n1006_));
  NAND2_X1  g0878(.A1(new_n1004_), .A2(new_n1006_), .ZN(new_n1007_));
  NAND3_X1  g0879(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n1008_));
  NOR2_X1   g0880(.A1(new_n853_), .A2(new_n849_), .ZN(new_n1009_));
  NAND2_X1  g0881(.A1(new_n773_), .A2(new_n1009_), .ZN(new_n1010_));
  NAND2_X1  g0882(.A1(new_n1008_), .A2(new_n1010_), .ZN(new_n1011_));
  AOI22_X1  g0883(.A1(new_n997_), .A2(new_n998_), .B1(new_n1001_), .B2(new_n1002_), .ZN(new_n1012_));
  NAND3_X1  g0884(.A1(new_n1012_), .A2(new_n1005_), .A3(new_n1000_), .ZN(new_n1013_));
  NAND3_X1  g0885(.A1(new_n1007_), .A2(new_n1011_), .A3(new_n1013_), .ZN(new_n1014_));
  INV_X1    g0886(.A(new_n1014_), .ZN(new_n1015_));
  AOI21_X1  g0887(.A(new_n1011_), .B1(new_n1007_), .B2(new_n1013_), .ZN(new_n1016_));
  OAI21_X1  g0888(.A(new_n896_), .B1(new_n1015_), .B2(new_n1016_), .ZN(new_n1017_));
  INV_X1    g0889(.A(new_n1011_), .ZN(new_n1018_));
  NOR2_X1   g0890(.A1(new_n1004_), .A2(new_n1006_), .ZN(new_n1019_));
  AOI21_X1  g0891(.A(new_n1005_), .B1(new_n1012_), .B2(new_n1000_), .ZN(new_n1020_));
  OAI21_X1  g0892(.A(new_n1018_), .B1(new_n1019_), .B2(new_n1020_), .ZN(new_n1021_));
  INV_X1    g0893(.A(new_n896_), .ZN(new_n1022_));
  NAND3_X1  g0894(.A1(new_n1021_), .A2(new_n1022_), .A3(new_n1014_), .ZN(new_n1023_));
  NAND2_X1  g0895(.A1(new_n1017_), .A2(new_n1023_), .ZN(new_n1024_));
  OAI21_X1  g0896(.A(new_n859_), .B1(new_n867_), .B2(new_n861_), .ZN(new_n1025_));
  INV_X1    g0897(.A(new_n1025_), .ZN(new_n1026_));
  NAND2_X1  g0898(.A1(new_n1024_), .A2(new_n1026_), .ZN(new_n1027_));
  NOR2_X1   g0899(.A1(new_n165_), .A2(new_n648_), .ZN(new_n1028_));
  INV_X1    g0900(.A(new_n1028_), .ZN(new_n1029_));
  NAND3_X1  g0901(.A1(new_n1017_), .A2(new_n1023_), .A3(new_n1025_), .ZN(new_n1030_));
  NAND3_X1  g0902(.A1(new_n1027_), .A2(new_n1029_), .A3(new_n1030_), .ZN(new_n1031_));
  AND3_X1   g0903(.A1(new_n1017_), .A2(new_n1023_), .A3(new_n1025_), .ZN(new_n1032_));
  AOI21_X1  g0904(.A(new_n1025_), .B1(new_n1017_), .B2(new_n1023_), .ZN(new_n1033_));
  OAI21_X1  g0905(.A(new_n1028_), .B1(new_n1032_), .B2(new_n1033_), .ZN(new_n1034_));
  NAND3_X1  g0906(.A1(new_n895_), .A2(new_n1031_), .A3(new_n1034_), .ZN(new_n1035_));
  NAND2_X1  g0907(.A1(new_n873_), .A2(new_n871_), .ZN(new_n1036_));
  INV_X1    g0908(.A(new_n1036_), .ZN(new_n1037_));
  NAND2_X1  g0909(.A1(new_n1035_), .A2(new_n1037_), .ZN(new_n1038_));
  NOR2_X1   g0910(.A1(new_n218_), .A2(new_n654_), .ZN(new_n1039_));
  INV_X1    g0911(.A(new_n1039_), .ZN(new_n1040_));
  NAND4_X1  g0912(.A1(new_n1036_), .A2(new_n895_), .A3(new_n1031_), .A4(new_n1034_), .ZN(new_n1041_));
  NAND3_X1  g0913(.A1(new_n1038_), .A2(new_n1040_), .A3(new_n1041_), .ZN(new_n1042_));
  NAND2_X1  g0914(.A1(new_n1038_), .A2(new_n1041_), .ZN(new_n1043_));
  NAND2_X1  g0915(.A1(new_n1043_), .A2(new_n1039_), .ZN(new_n1044_));
  NAND3_X1  g0916(.A1(new_n894_), .A2(new_n1042_), .A3(new_n1044_), .ZN(new_n1045_));
  INV_X1    g0917(.A(new_n1045_), .ZN(new_n1046_));
  AOI21_X1  g0918(.A(new_n894_), .B1(new_n1042_), .B2(new_n1044_), .ZN(new_n1047_));
  NOR2_X1   g0919(.A1(new_n1046_), .A2(new_n1047_), .ZN(new_n1048_));
  NOR2_X1   g0920(.A1(new_n132_), .A2(new_n890_), .ZN(new_n1049_));
  INV_X1    g0921(.A(new_n1049_), .ZN(new_n1050_));
  NAND2_X1  g0922(.A1(new_n1048_), .A2(new_n1050_), .ZN(new_n1051_));
  OAI21_X1  g0923(.A(new_n1049_), .B1(new_n1046_), .B2(new_n1047_), .ZN(new_n1052_));
  NAND3_X1  g0924(.A1(new_n893_), .A2(new_n1051_), .A3(new_n1052_), .ZN(new_n1053_));
  INV_X1    g0925(.A(new_n1053_), .ZN(new_n1054_));
  AOI21_X1  g0926(.A(new_n893_), .B1(new_n1052_), .B2(new_n1051_), .ZN(new_n1055_));
  NOR2_X1   g0927(.A1(new_n1054_), .A2(new_n1055_), .ZN(new_n1056_));
  INV_X1    g0928(.A(G494gat), .ZN(new_n1057_));
  NOR2_X1   g0929(.A1(new_n129_), .A2(new_n1057_), .ZN(new_n1058_));
  INV_X1    g0930(.A(new_n1058_), .ZN(new_n1059_));
  XNOR2_X1  g0931(.A(new_n1056_), .B(new_n1059_), .ZN(G5672gat));
  OAI21_X1  g0932(.A(new_n1053_), .B1(new_n1055_), .B2(new_n1058_), .ZN(new_n1061_));
  OAI21_X1  g0933(.A(new_n1045_), .B1(new_n1047_), .B2(new_n1049_), .ZN(new_n1062_));
  NAND3_X1  g0934(.A1(new_n1036_), .A2(new_n1031_), .A3(new_n1034_), .ZN(new_n1063_));
  NAND2_X1  g0935(.A1(new_n1042_), .A2(new_n1063_), .ZN(new_n1064_));
  NOR2_X1   g0936(.A1(new_n166_), .A2(new_n648_), .ZN(new_n1065_));
  NOR2_X1   g0937(.A1(new_n242_), .A2(new_n533_), .ZN(new_n1066_));
  NOR2_X1   g0938(.A1(new_n243_), .A2(new_n443_), .ZN(new_n1067_));
  NOR2_X1   g0939(.A1(new_n300_), .A2(new_n363_), .ZN(new_n1068_));
  NAND2_X1  g0940(.A1(new_n950_), .A2(new_n948_), .ZN(new_n1069_));
  NAND2_X1  g0941(.A1(G222gat), .A2(G290gat), .ZN(new_n1070_));
  NAND2_X1  g0942(.A1(G239gat), .A2(G273gat), .ZN(new_n1071_));
  NAND2_X1  g0943(.A1(new_n1070_), .A2(new_n1071_), .ZN(new_n1072_));
  NAND4_X1  g0944(.A1(G222gat), .A2(G239gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1073_));
  NAND2_X1  g0945(.A1(new_n1072_), .A2(new_n1073_), .ZN(new_n1074_));
  NAND2_X1  g0946(.A1(new_n1074_), .A2(new_n907_), .ZN(new_n1075_));
  NAND2_X1  g0947(.A1(new_n908_), .A2(new_n1073_), .ZN(new_n1076_));
  NAND2_X1  g0948(.A1(new_n1075_), .A2(new_n1076_), .ZN(new_n1077_));
  NAND2_X1  g0949(.A1(G205gat), .A2(G307gat), .ZN(new_n1078_));
  INV_X1    g0950(.A(new_n1078_), .ZN(new_n1079_));
  NAND2_X1  g0951(.A1(new_n1077_), .A2(new_n1079_), .ZN(new_n1080_));
  NAND3_X1  g0952(.A1(new_n1075_), .A2(new_n1078_), .A3(new_n1076_), .ZN(new_n1081_));
  NAND2_X1  g0953(.A1(new_n1080_), .A2(new_n1081_), .ZN(new_n1082_));
  NAND3_X1  g0954(.A1(new_n1082_), .A2(new_n906_), .A3(new_n916_), .ZN(new_n1083_));
  INV_X1    g0955(.A(G188gat), .ZN(new_n1084_));
  NOR2_X1   g0956(.A1(new_n1084_), .A2(new_n159_), .ZN(new_n1085_));
  INV_X1    g0957(.A(new_n1085_), .ZN(new_n1086_));
  INV_X1    g0958(.A(new_n906_), .ZN(new_n1087_));
  NAND3_X1  g0959(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n1088_));
  AOI21_X1  g0960(.A(new_n1087_), .B1(new_n1088_), .B2(new_n911_), .ZN(new_n1089_));
  OAI211_X1 g0961(.A(new_n1083_), .B(new_n1086_), .C1(new_n1082_), .C2(new_n1089_), .ZN(new_n1090_));
  INV_X1    g0962(.A(new_n1090_), .ZN(new_n1091_));
  OR2_X1    g0963(.A1(new_n1089_), .A2(new_n1082_), .ZN(new_n1092_));
  AOI21_X1  g0964(.A(new_n1086_), .B1(new_n1092_), .B2(new_n1083_), .ZN(new_n1093_));
  NOR2_X1   g0965(.A1(new_n1091_), .A2(new_n1093_), .ZN(new_n1094_));
  NOR2_X1   g0966(.A1(new_n926_), .A2(new_n915_), .ZN(new_n1095_));
  INV_X1    g0967(.A(new_n1095_), .ZN(new_n1096_));
  AOI21_X1  g0968(.A(KEYINPUT33), .B1(new_n933_), .B2(new_n1096_), .ZN(new_n1097_));
  INV_X1    g0969(.A(KEYINPUT33), .ZN(new_n1098_));
  AOI211_X1 g0970(.A(new_n1098_), .B(new_n1095_), .C1(new_n930_), .C2(new_n932_), .ZN(new_n1099_));
  OAI21_X1  g0971(.A(new_n1094_), .B1(new_n1097_), .B2(new_n1099_), .ZN(new_n1100_));
  NOR2_X1   g0972(.A1(new_n543_), .A2(new_n198_), .ZN(new_n1101_));
  AOI21_X1  g0973(.A(new_n1095_), .B1(new_n930_), .B2(new_n932_), .ZN(new_n1102_));
  NAND2_X1  g0974(.A1(new_n1102_), .A2(KEYINPUT33), .ZN(new_n1103_));
  OR2_X1    g0975(.A1(new_n1091_), .A2(new_n1093_), .ZN(new_n1104_));
  NAND2_X1  g0976(.A1(new_n1103_), .A2(new_n1104_), .ZN(new_n1105_));
  AND3_X1   g0977(.A1(new_n1100_), .A2(new_n1101_), .A3(new_n1105_), .ZN(new_n1106_));
  AOI21_X1  g0978(.A(new_n1101_), .B1(new_n1100_), .B2(new_n1105_), .ZN(new_n1107_));
  OAI21_X1  g0979(.A(new_n1069_), .B1(new_n1106_), .B2(new_n1107_), .ZN(new_n1108_));
  INV_X1    g0980(.A(new_n1101_), .ZN(new_n1109_));
  INV_X1    g0981(.A(new_n917_), .ZN(new_n1110_));
  AOI21_X1  g0982(.A(new_n1110_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n1111_));
  OAI21_X1  g0983(.A(new_n1096_), .B1(new_n1111_), .B2(new_n931_), .ZN(new_n1112_));
  NAND2_X1  g0984(.A1(new_n1112_), .A2(new_n1098_), .ZN(new_n1113_));
  AOI21_X1  g0985(.A(new_n1104_), .B1(new_n1113_), .B2(new_n1103_), .ZN(new_n1114_));
  NOR2_X1   g0986(.A1(new_n1099_), .A2(new_n1094_), .ZN(new_n1115_));
  OAI21_X1  g0987(.A(new_n1109_), .B1(new_n1114_), .B2(new_n1115_), .ZN(new_n1116_));
  NAND3_X1  g0988(.A1(new_n1100_), .A2(new_n1101_), .A3(new_n1105_), .ZN(new_n1117_));
  NAND4_X1  g0989(.A1(new_n1116_), .A2(new_n948_), .A3(new_n953_), .A4(new_n1117_), .ZN(new_n1118_));
  NAND2_X1  g0990(.A1(new_n1108_), .A2(new_n1118_), .ZN(new_n1119_));
  NOR2_X1   g0991(.A1(new_n542_), .A2(new_n276_), .ZN(new_n1120_));
  INV_X1    g0992(.A(new_n1120_), .ZN(new_n1121_));
  NAND2_X1  g0993(.A1(new_n1119_), .A2(new_n1121_), .ZN(new_n1122_));
  NAND3_X1  g0994(.A1(new_n1108_), .A2(new_n1118_), .A3(new_n1120_), .ZN(new_n1123_));
  NAND3_X1  g0995(.A1(new_n938_), .A2(new_n939_), .A3(new_n953_), .ZN(new_n1124_));
  AND3_X1   g0996(.A1(new_n962_), .A2(KEYINPUT34), .A3(new_n1124_), .ZN(new_n1125_));
  AOI21_X1  g0997(.A(KEYINPUT34), .B1(new_n962_), .B2(new_n1124_), .ZN(new_n1126_));
  OAI211_X1 g0998(.A(new_n1122_), .B(new_n1123_), .C1(new_n1125_), .C2(new_n1126_), .ZN(new_n1127_));
  AND3_X1   g0999(.A1(new_n1108_), .A2(new_n1118_), .A3(new_n1120_), .ZN(new_n1128_));
  AOI21_X1  g1000(.A(new_n1120_), .B1(new_n1108_), .B2(new_n1118_), .ZN(new_n1129_));
  INV_X1    g1001(.A(KEYINPUT34), .ZN(new_n1130_));
  NAND2_X1  g1002(.A1(new_n962_), .A2(new_n1124_), .ZN(new_n1131_));
  OAI22_X1  g1003(.A1(new_n1128_), .A2(new_n1129_), .B1(new_n1130_), .B2(new_n1131_), .ZN(new_n1132_));
  NOR2_X1   g1004(.A1(new_n377_), .A2(new_n289_), .ZN(new_n1133_));
  AND3_X1   g1005(.A1(new_n1127_), .A2(new_n1132_), .A3(new_n1133_), .ZN(new_n1134_));
  AOI21_X1  g1006(.A(new_n1133_), .B1(new_n1127_), .B2(new_n1132_), .ZN(new_n1135_));
  NAND2_X1  g1007(.A1(new_n980_), .A2(new_n979_), .ZN(new_n1136_));
  INV_X1    g1008(.A(new_n1136_), .ZN(new_n1137_));
  NOR3_X1   g1009(.A1(new_n1134_), .A2(new_n1135_), .A3(new_n1137_), .ZN(new_n1138_));
  NAND2_X1  g1010(.A1(new_n1127_), .A2(new_n1132_), .ZN(new_n1139_));
  INV_X1    g1011(.A(new_n1133_), .ZN(new_n1140_));
  NAND2_X1  g1012(.A1(new_n1139_), .A2(new_n1140_), .ZN(new_n1141_));
  NAND3_X1  g1013(.A1(new_n1127_), .A2(new_n1133_), .A3(new_n1132_), .ZN(new_n1142_));
  AOI21_X1  g1014(.A(new_n1136_), .B1(new_n1141_), .B2(new_n1142_), .ZN(new_n1143_));
  OAI21_X1  g1015(.A(new_n1068_), .B1(new_n1138_), .B2(new_n1143_), .ZN(new_n1144_));
  NAND2_X1  g1016(.A1(new_n971_), .A2(new_n980_), .ZN(new_n1145_));
  OR2_X1    g1017(.A1(new_n1145_), .A2(KEYINPUT32), .ZN(new_n1146_));
  NAND2_X1  g1018(.A1(new_n1145_), .A2(KEYINPUT32), .ZN(new_n1147_));
  NAND3_X1  g1019(.A1(new_n1146_), .A2(new_n986_), .A3(new_n1147_), .ZN(new_n1148_));
  NAND3_X1  g1020(.A1(new_n984_), .A2(new_n987_), .A3(new_n991_), .ZN(new_n1149_));
  NAND2_X1  g1021(.A1(new_n1148_), .A2(new_n1149_), .ZN(new_n1150_));
  OAI21_X1  g1022(.A(new_n1137_), .B1(new_n1134_), .B2(new_n1135_), .ZN(new_n1151_));
  NAND3_X1  g1023(.A1(new_n1141_), .A2(new_n1136_), .A3(new_n1142_), .ZN(new_n1152_));
  INV_X1    g1024(.A(new_n1068_), .ZN(new_n1153_));
  NAND3_X1  g1025(.A1(new_n1151_), .A2(new_n1152_), .A3(new_n1153_), .ZN(new_n1154_));
  AND3_X1   g1026(.A1(new_n1144_), .A2(new_n1150_), .A3(new_n1154_), .ZN(new_n1155_));
  AOI21_X1  g1027(.A(new_n1150_), .B1(new_n1144_), .B2(new_n1154_), .ZN(new_n1156_));
  OAI21_X1  g1028(.A(new_n1067_), .B1(new_n1155_), .B2(new_n1156_), .ZN(new_n1157_));
  NAND2_X1  g1029(.A1(new_n1144_), .A2(new_n1154_), .ZN(new_n1158_));
  INV_X1    g1030(.A(new_n1150_), .ZN(new_n1159_));
  NAND2_X1  g1031(.A1(new_n1158_), .A2(new_n1159_), .ZN(new_n1160_));
  INV_X1    g1032(.A(new_n1067_), .ZN(new_n1161_));
  NAND3_X1  g1033(.A1(new_n1144_), .A2(new_n1150_), .A3(new_n1154_), .ZN(new_n1162_));
  NAND3_X1  g1034(.A1(new_n1160_), .A2(new_n1161_), .A3(new_n1162_), .ZN(new_n1163_));
  NAND2_X1  g1035(.A1(new_n1157_), .A2(new_n1163_), .ZN(new_n1164_));
  XOR2_X1   g1036(.A(new_n1002_), .B(KEYINPUT31), .Z(new_n1165_));
  OR2_X1    g1037(.A1(new_n1165_), .A2(new_n1001_), .ZN(new_n1166_));
  AND3_X1   g1038(.A1(new_n1007_), .A2(new_n1164_), .A3(new_n1166_), .ZN(new_n1167_));
  AOI21_X1  g1039(.A(new_n1164_), .B1(new_n1007_), .B2(new_n1166_), .ZN(new_n1168_));
  OAI21_X1  g1040(.A(new_n1066_), .B1(new_n1167_), .B2(new_n1168_), .ZN(new_n1169_));
  OAI21_X1  g1041(.A(new_n1014_), .B1(new_n1016_), .B2(new_n896_), .ZN(new_n1170_));
  NOR2_X1   g1042(.A1(new_n1165_), .A2(new_n1001_), .ZN(new_n1171_));
  OAI211_X1 g1043(.A(new_n1163_), .B(new_n1157_), .C1(new_n1020_), .C2(new_n1171_), .ZN(new_n1172_));
  INV_X1    g1044(.A(new_n1066_), .ZN(new_n1173_));
  NAND3_X1  g1045(.A1(new_n1007_), .A2(new_n1164_), .A3(new_n1166_), .ZN(new_n1174_));
  NAND3_X1  g1046(.A1(new_n1172_), .A2(new_n1173_), .A3(new_n1174_), .ZN(new_n1175_));
  AND3_X1   g1047(.A1(new_n1169_), .A2(new_n1170_), .A3(new_n1175_), .ZN(new_n1176_));
  AOI21_X1  g1048(.A(new_n1170_), .B1(new_n1169_), .B2(new_n1175_), .ZN(new_n1177_));
  OAI21_X1  g1049(.A(new_n1065_), .B1(new_n1176_), .B2(new_n1177_), .ZN(new_n1178_));
  OAI21_X1  g1050(.A(new_n1030_), .B1(new_n1033_), .B2(new_n1028_), .ZN(new_n1179_));
  INV_X1    g1051(.A(new_n1170_), .ZN(new_n1180_));
  NOR3_X1   g1052(.A1(new_n1167_), .A2(new_n1168_), .A3(new_n1066_), .ZN(new_n1181_));
  AOI21_X1  g1053(.A(new_n1173_), .B1(new_n1172_), .B2(new_n1174_), .ZN(new_n1182_));
  OAI21_X1  g1054(.A(new_n1180_), .B1(new_n1181_), .B2(new_n1182_), .ZN(new_n1183_));
  INV_X1    g1055(.A(new_n1065_), .ZN(new_n1184_));
  NAND3_X1  g1056(.A1(new_n1169_), .A2(new_n1170_), .A3(new_n1175_), .ZN(new_n1185_));
  NAND3_X1  g1057(.A1(new_n1183_), .A2(new_n1184_), .A3(new_n1185_), .ZN(new_n1186_));
  AND3_X1   g1058(.A1(new_n1178_), .A2(new_n1179_), .A3(new_n1186_), .ZN(new_n1187_));
  AOI21_X1  g1059(.A(new_n1179_), .B1(new_n1178_), .B2(new_n1186_), .ZN(new_n1188_));
  NOR2_X1   g1060(.A1(new_n165_), .A2(new_n654_), .ZN(new_n1189_));
  NOR3_X1   g1061(.A1(new_n1187_), .A2(new_n1188_), .A3(new_n1189_), .ZN(new_n1190_));
  INV_X1    g1062(.A(new_n1189_), .ZN(new_n1191_));
  AOI21_X1  g1063(.A(new_n1032_), .B1(new_n1027_), .B2(new_n1029_), .ZN(new_n1192_));
  NOR3_X1   g1064(.A1(new_n1176_), .A2(new_n1177_), .A3(new_n1065_), .ZN(new_n1193_));
  AOI21_X1  g1065(.A(new_n1184_), .B1(new_n1183_), .B2(new_n1185_), .ZN(new_n1194_));
  OAI21_X1  g1066(.A(new_n1192_), .B1(new_n1193_), .B2(new_n1194_), .ZN(new_n1195_));
  NAND3_X1  g1067(.A1(new_n1178_), .A2(new_n1179_), .A3(new_n1186_), .ZN(new_n1196_));
  AOI21_X1  g1068(.A(new_n1191_), .B1(new_n1195_), .B2(new_n1196_), .ZN(new_n1197_));
  NOR2_X1   g1069(.A1(new_n1190_), .A2(new_n1197_), .ZN(new_n1198_));
  NAND2_X1  g1070(.A1(new_n1064_), .A2(new_n1198_), .ZN(new_n1199_));
  NOR2_X1   g1071(.A1(new_n218_), .A2(new_n890_), .ZN(new_n1200_));
  INV_X1    g1072(.A(new_n1200_), .ZN(new_n1201_));
  OAI211_X1 g1073(.A(new_n1042_), .B(new_n1063_), .C1(new_n1190_), .C2(new_n1197_), .ZN(new_n1202_));
  NAND3_X1  g1074(.A1(new_n1199_), .A2(new_n1201_), .A3(new_n1202_), .ZN(new_n1203_));
  INV_X1    g1075(.A(new_n1199_), .ZN(new_n1204_));
  INV_X1    g1076(.A(new_n1202_), .ZN(new_n1205_));
  OAI21_X1  g1077(.A(new_n1200_), .B1(new_n1204_), .B2(new_n1205_), .ZN(new_n1206_));
  AOI21_X1  g1078(.A(new_n1062_), .B1(new_n1203_), .B2(new_n1206_), .ZN(new_n1207_));
  INV_X1    g1079(.A(new_n1207_), .ZN(new_n1208_));
  NAND3_X1  g1080(.A1(new_n1062_), .A2(new_n1206_), .A3(new_n1203_), .ZN(new_n1209_));
  OAI211_X1 g1081(.A(new_n1208_), .B(new_n1209_), .C1(new_n132_), .C2(new_n1057_), .ZN(new_n1210_));
  NOR2_X1   g1082(.A1(new_n132_), .A2(new_n1057_), .ZN(new_n1211_));
  INV_X1    g1083(.A(new_n1209_), .ZN(new_n1212_));
  OAI21_X1  g1084(.A(new_n1211_), .B1(new_n1212_), .B2(new_n1207_), .ZN(new_n1213_));
  AOI21_X1  g1085(.A(new_n1061_), .B1(new_n1210_), .B2(new_n1213_), .ZN(new_n1214_));
  INV_X1    g1086(.A(new_n1214_), .ZN(new_n1215_));
  NAND3_X1  g1087(.A1(new_n1061_), .A2(new_n1213_), .A3(new_n1210_), .ZN(new_n1216_));
  NAND2_X1  g1088(.A1(new_n1215_), .A2(new_n1216_), .ZN(new_n1217_));
  INV_X1    g1089(.A(G511gat), .ZN(new_n1218_));
  NOR2_X1   g1090(.A1(new_n129_), .A2(new_n1218_), .ZN(new_n1219_));
  XNOR2_X1  g1091(.A(new_n1217_), .B(new_n1219_), .ZN(G5971gat));
  OAI21_X1  g1092(.A(new_n1216_), .B1(new_n1214_), .B2(new_n1219_), .ZN(new_n1221_));
  OAI21_X1  g1093(.A(new_n1209_), .B1(new_n1207_), .B2(new_n1211_), .ZN(new_n1222_));
  OAI21_X1  g1094(.A(new_n1199_), .B1(new_n1205_), .B2(new_n1200_), .ZN(new_n1223_));
  NAND2_X1  g1095(.A1(G52gat), .A2(G477gat), .ZN(new_n1224_));
  XNOR2_X1  g1096(.A(new_n1224_), .B(KEYINPUT39), .ZN(new_n1225_));
  INV_X1    g1097(.A(new_n1225_), .ZN(new_n1226_));
  AOI21_X1  g1098(.A(new_n1187_), .B1(new_n1191_), .B2(new_n1195_), .ZN(new_n1227_));
  AOI21_X1  g1099(.A(new_n1176_), .B1(new_n1184_), .B2(new_n1183_), .ZN(new_n1228_));
  AOI21_X1  g1100(.A(new_n1168_), .B1(new_n1174_), .B2(new_n1173_), .ZN(new_n1229_));
  AOI21_X1  g1101(.A(new_n1155_), .B1(new_n1160_), .B2(new_n1161_), .ZN(new_n1230_));
  NAND3_X1  g1102(.A1(new_n1116_), .A2(new_n1117_), .A3(new_n1069_), .ZN(new_n1231_));
  INV_X1    g1103(.A(G256gat), .ZN(new_n1232_));
  NOR2_X1   g1104(.A1(new_n1073_), .A2(new_n1232_), .ZN(new_n1233_));
  INV_X1    g1105(.A(new_n1233_), .ZN(new_n1234_));
  NAND2_X1  g1106(.A1(new_n1234_), .A2(KEYINPUT37), .ZN(new_n1235_));
  NAND2_X1  g1107(.A1(G239gat), .A2(G290gat), .ZN(new_n1236_));
  NAND3_X1  g1108(.A1(new_n1236_), .A2(G256gat), .A3(G273gat), .ZN(new_n1237_));
  NAND2_X1  g1109(.A1(G256gat), .A2(G273gat), .ZN(new_n1238_));
  NAND3_X1  g1110(.A1(new_n1238_), .A2(G239gat), .A3(G290gat), .ZN(new_n1239_));
  NAND2_X1  g1111(.A1(new_n1237_), .A2(new_n1239_), .ZN(new_n1240_));
  AOI21_X1  g1112(.A(new_n1233_), .B1(new_n1240_), .B2(new_n1073_), .ZN(new_n1241_));
  OAI21_X1  g1113(.A(new_n1235_), .B1(new_n1241_), .B2(KEYINPUT37), .ZN(new_n1242_));
  NAND2_X1  g1114(.A1(G222gat), .A2(G307gat), .ZN(new_n1243_));
  INV_X1    g1115(.A(new_n1243_), .ZN(new_n1244_));
  NAND2_X1  g1116(.A1(new_n1242_), .A2(new_n1244_), .ZN(new_n1245_));
  NAND2_X1  g1117(.A1(new_n1081_), .A2(new_n1075_), .ZN(new_n1246_));
  NAND2_X1  g1118(.A1(new_n1241_), .A2(new_n1243_), .ZN(new_n1247_));
  NAND3_X1  g1119(.A1(new_n1245_), .A2(new_n1246_), .A3(new_n1247_), .ZN(new_n1248_));
  NAND3_X1  g1120(.A1(new_n1074_), .A2(KEYINPUT36), .A3(new_n907_), .ZN(new_n1249_));
  INV_X1    g1121(.A(KEYINPUT36), .ZN(new_n1250_));
  NAND2_X1  g1122(.A1(new_n1075_), .A2(new_n1250_), .ZN(new_n1251_));
  AND3_X1   g1123(.A1(new_n1081_), .A2(new_n1249_), .A3(new_n1251_), .ZN(new_n1252_));
  XNOR2_X1  g1124(.A(new_n1236_), .B(new_n1238_), .ZN(new_n1253_));
  INV_X1    g1125(.A(new_n1073_), .ZN(new_n1254_));
  OAI21_X1  g1126(.A(new_n1234_), .B1(new_n1253_), .B2(new_n1254_), .ZN(new_n1255_));
  NAND2_X1  g1127(.A1(new_n1255_), .A2(new_n1243_), .ZN(new_n1256_));
  NAND2_X1  g1128(.A1(new_n1241_), .A2(new_n1244_), .ZN(new_n1257_));
  NAND3_X1  g1129(.A1(new_n1252_), .A2(new_n1256_), .A3(new_n1257_), .ZN(new_n1258_));
  NAND2_X1  g1130(.A1(new_n1248_), .A2(new_n1258_), .ZN(new_n1259_));
  INV_X1    g1131(.A(G205gat), .ZN(new_n1260_));
  NOR2_X1   g1132(.A1(new_n1260_), .A2(new_n159_), .ZN(new_n1261_));
  INV_X1    g1133(.A(new_n1261_), .ZN(new_n1262_));
  NAND2_X1  g1134(.A1(new_n1259_), .A2(new_n1262_), .ZN(new_n1263_));
  AND3_X1   g1135(.A1(new_n1082_), .A2(new_n906_), .A3(new_n916_), .ZN(new_n1264_));
  OAI21_X1  g1136(.A(new_n1092_), .B1(new_n1264_), .B2(new_n1085_), .ZN(new_n1265_));
  NAND3_X1  g1137(.A1(new_n1248_), .A2(new_n1258_), .A3(new_n1261_), .ZN(new_n1266_));
  NAND3_X1  g1138(.A1(new_n1263_), .A2(new_n1265_), .A3(new_n1266_), .ZN(new_n1267_));
  INV_X1    g1139(.A(new_n1267_), .ZN(new_n1268_));
  AOI21_X1  g1140(.A(new_n1265_), .B1(new_n1263_), .B2(new_n1266_), .ZN(new_n1269_));
  OAI22_X1  g1141(.A1(new_n1268_), .A2(new_n1269_), .B1(new_n1084_), .B2(new_n198_), .ZN(new_n1270_));
  INV_X1    g1142(.A(new_n1266_), .ZN(new_n1271_));
  AOI21_X1  g1143(.A(new_n1261_), .B1(new_n1248_), .B2(new_n1258_), .ZN(new_n1272_));
  OAI211_X1 g1144(.A(new_n1092_), .B(new_n1090_), .C1(new_n1271_), .C2(new_n1272_), .ZN(new_n1273_));
  NOR2_X1   g1145(.A1(new_n1084_), .A2(new_n198_), .ZN(new_n1274_));
  NAND3_X1  g1146(.A1(new_n1273_), .A2(new_n1274_), .A3(new_n1267_), .ZN(new_n1275_));
  NOR2_X1   g1147(.A1(new_n1104_), .A2(new_n1102_), .ZN(new_n1276_));
  OAI211_X1 g1148(.A(new_n1270_), .B(new_n1275_), .C1(new_n1107_), .C2(new_n1276_), .ZN(new_n1277_));
  INV_X1    g1149(.A(new_n1276_), .ZN(new_n1278_));
  INV_X1    g1150(.A(KEYINPUT38), .ZN(new_n1279_));
  NAND3_X1  g1151(.A1(new_n1270_), .A2(new_n1275_), .A3(new_n1279_), .ZN(new_n1280_));
  OAI221_X1 g1152(.A(KEYINPUT38), .B1(new_n1084_), .B2(new_n198_), .C1(new_n1268_), .C2(new_n1269_), .ZN(new_n1281_));
  NAND4_X1  g1153(.A1(new_n1116_), .A2(new_n1278_), .A3(new_n1280_), .A4(new_n1281_), .ZN(new_n1282_));
  NOR2_X1   g1154(.A1(new_n543_), .A2(new_n276_), .ZN(new_n1283_));
  NAND3_X1  g1155(.A1(new_n1277_), .A2(new_n1282_), .A3(new_n1283_), .ZN(new_n1284_));
  INV_X1    g1156(.A(new_n1284_), .ZN(new_n1285_));
  AOI21_X1  g1157(.A(new_n1283_), .B1(new_n1277_), .B2(new_n1282_), .ZN(new_n1286_));
  OAI211_X1 g1158(.A(new_n1122_), .B(new_n1231_), .C1(new_n1285_), .C2(new_n1286_), .ZN(new_n1287_));
  NAND2_X1  g1159(.A1(new_n1277_), .A2(new_n1282_), .ZN(new_n1288_));
  INV_X1    g1160(.A(new_n1283_), .ZN(new_n1289_));
  NAND2_X1  g1161(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_));
  INV_X1    g1162(.A(new_n1231_), .ZN(new_n1291_));
  OAI211_X1 g1163(.A(new_n1290_), .B(new_n1284_), .C1(new_n1129_), .C2(new_n1291_), .ZN(new_n1292_));
  NAND2_X1  g1164(.A1(new_n1287_), .A2(new_n1292_), .ZN(new_n1293_));
  NOR2_X1   g1165(.A1(new_n542_), .A2(new_n289_), .ZN(new_n1294_));
  NAND2_X1  g1166(.A1(new_n1293_), .A2(new_n1294_), .ZN(new_n1295_));
  INV_X1    g1167(.A(new_n1294_), .ZN(new_n1296_));
  NAND3_X1  g1168(.A1(new_n1287_), .A2(new_n1292_), .A3(new_n1296_), .ZN(new_n1297_));
  NAND3_X1  g1169(.A1(new_n1122_), .A2(new_n1123_), .A3(new_n1131_), .ZN(new_n1298_));
  INV_X1    g1170(.A(new_n1298_), .ZN(new_n1299_));
  OAI211_X1 g1171(.A(new_n1295_), .B(new_n1297_), .C1(new_n1135_), .C2(new_n1299_), .ZN(new_n1300_));
  AND3_X1   g1172(.A1(new_n1287_), .A2(new_n1292_), .A3(new_n1296_), .ZN(new_n1301_));
  AOI21_X1  g1173(.A(new_n1296_), .B1(new_n1287_), .B2(new_n1292_), .ZN(new_n1302_));
  OAI211_X1 g1174(.A(new_n1141_), .B(new_n1298_), .C1(new_n1301_), .C2(new_n1302_), .ZN(new_n1303_));
  NAND2_X1  g1175(.A1(new_n1300_), .A2(new_n1303_), .ZN(new_n1304_));
  NOR2_X1   g1176(.A1(new_n377_), .A2(new_n363_), .ZN(new_n1305_));
  NAND2_X1  g1177(.A1(new_n1304_), .A2(new_n1305_), .ZN(new_n1306_));
  NAND2_X1  g1178(.A1(new_n1154_), .A2(KEYINPUT35), .ZN(new_n1307_));
  INV_X1    g1179(.A(new_n1305_), .ZN(new_n1308_));
  NAND3_X1  g1180(.A1(new_n1300_), .A2(new_n1303_), .A3(new_n1308_), .ZN(new_n1309_));
  NAND3_X1  g1181(.A1(new_n1306_), .A2(new_n1307_), .A3(new_n1309_), .ZN(new_n1310_));
  NAND2_X1  g1182(.A1(new_n1154_), .A2(new_n1152_), .ZN(new_n1311_));
  INV_X1    g1183(.A(new_n1311_), .ZN(new_n1312_));
  NAND2_X1  g1184(.A1(new_n1310_), .A2(new_n1312_), .ZN(new_n1313_));
  NOR2_X1   g1185(.A1(new_n300_), .A2(new_n443_), .ZN(new_n1314_));
  INV_X1    g1186(.A(new_n1314_), .ZN(new_n1315_));
  NAND4_X1  g1187(.A1(new_n1306_), .A2(new_n1311_), .A3(new_n1307_), .A4(new_n1309_), .ZN(new_n1316_));
  AND3_X1   g1188(.A1(new_n1313_), .A2(new_n1315_), .A3(new_n1316_), .ZN(new_n1317_));
  AOI21_X1  g1189(.A(new_n1315_), .B1(new_n1313_), .B2(new_n1316_), .ZN(new_n1318_));
  OAI21_X1  g1190(.A(new_n1230_), .B1(new_n1317_), .B2(new_n1318_), .ZN(new_n1319_));
  NOR2_X1   g1191(.A1(new_n243_), .A2(new_n533_), .ZN(new_n1320_));
  INV_X1    g1192(.A(new_n1320_), .ZN(new_n1321_));
  AND3_X1   g1193(.A1(new_n1300_), .A2(new_n1303_), .A3(new_n1308_), .ZN(new_n1322_));
  AOI21_X1  g1194(.A(new_n1308_), .B1(new_n1300_), .B2(new_n1303_), .ZN(new_n1323_));
  NOR2_X1   g1195(.A1(new_n1322_), .A2(new_n1323_), .ZN(new_n1324_));
  AOI21_X1  g1196(.A(new_n1311_), .B1(new_n1324_), .B2(new_n1307_), .ZN(new_n1325_));
  AND4_X1   g1197(.A1(new_n1311_), .A2(new_n1306_), .A3(new_n1307_), .A4(new_n1309_), .ZN(new_n1326_));
  OAI21_X1  g1198(.A(new_n1314_), .B1(new_n1325_), .B2(new_n1326_), .ZN(new_n1327_));
  INV_X1    g1199(.A(new_n1230_), .ZN(new_n1328_));
  NAND3_X1  g1200(.A1(new_n1313_), .A2(new_n1315_), .A3(new_n1316_), .ZN(new_n1329_));
  NAND3_X1  g1201(.A1(new_n1327_), .A2(new_n1328_), .A3(new_n1329_), .ZN(new_n1330_));
  AND3_X1   g1202(.A1(new_n1319_), .A2(new_n1321_), .A3(new_n1330_), .ZN(new_n1331_));
  AOI21_X1  g1203(.A(new_n1321_), .B1(new_n1319_), .B2(new_n1330_), .ZN(new_n1332_));
  OAI21_X1  g1204(.A(new_n1229_), .B1(new_n1331_), .B2(new_n1332_), .ZN(new_n1333_));
  NOR2_X1   g1205(.A1(new_n242_), .A2(new_n648_), .ZN(new_n1334_));
  INV_X1    g1206(.A(new_n1334_), .ZN(new_n1335_));
  OAI21_X1  g1207(.A(new_n1172_), .B1(new_n1167_), .B2(new_n1066_), .ZN(new_n1336_));
  NOR3_X1   g1208(.A1(new_n1317_), .A2(new_n1318_), .A3(new_n1230_), .ZN(new_n1337_));
  AOI21_X1  g1209(.A(new_n1328_), .B1(new_n1327_), .B2(new_n1329_), .ZN(new_n1338_));
  OAI21_X1  g1210(.A(new_n1320_), .B1(new_n1337_), .B2(new_n1338_), .ZN(new_n1339_));
  NAND3_X1  g1211(.A1(new_n1319_), .A2(new_n1321_), .A3(new_n1330_), .ZN(new_n1340_));
  NAND3_X1  g1212(.A1(new_n1336_), .A2(new_n1339_), .A3(new_n1340_), .ZN(new_n1341_));
  AND3_X1   g1213(.A1(new_n1333_), .A2(new_n1335_), .A3(new_n1341_), .ZN(new_n1342_));
  AOI21_X1  g1214(.A(new_n1335_), .B1(new_n1333_), .B2(new_n1341_), .ZN(new_n1343_));
  OAI21_X1  g1215(.A(new_n1228_), .B1(new_n1342_), .B2(new_n1343_), .ZN(new_n1344_));
  NOR2_X1   g1216(.A1(new_n166_), .A2(new_n654_), .ZN(new_n1345_));
  INV_X1    g1217(.A(new_n1345_), .ZN(new_n1346_));
  NAND2_X1  g1218(.A1(new_n1333_), .A2(new_n1341_), .ZN(new_n1347_));
  NAND2_X1  g1219(.A1(new_n1347_), .A2(new_n1334_), .ZN(new_n1348_));
  OAI21_X1  g1220(.A(new_n1185_), .B1(new_n1177_), .B2(new_n1065_), .ZN(new_n1349_));
  NAND3_X1  g1221(.A1(new_n1333_), .A2(new_n1341_), .A3(new_n1335_), .ZN(new_n1350_));
  NAND3_X1  g1222(.A1(new_n1348_), .A2(new_n1349_), .A3(new_n1350_), .ZN(new_n1351_));
  AND3_X1   g1223(.A1(new_n1344_), .A2(new_n1346_), .A3(new_n1351_), .ZN(new_n1352_));
  AOI21_X1  g1224(.A(new_n1346_), .B1(new_n1344_), .B2(new_n1351_), .ZN(new_n1353_));
  OAI21_X1  g1225(.A(new_n1227_), .B1(new_n1352_), .B2(new_n1353_), .ZN(new_n1354_));
  AND3_X1   g1226(.A1(new_n1348_), .A2(new_n1349_), .A3(new_n1350_), .ZN(new_n1355_));
  AOI21_X1  g1227(.A(new_n1349_), .B1(new_n1348_), .B2(new_n1350_), .ZN(new_n1356_));
  OAI21_X1  g1228(.A(new_n1345_), .B1(new_n1355_), .B2(new_n1356_), .ZN(new_n1357_));
  OAI21_X1  g1229(.A(new_n1196_), .B1(new_n1188_), .B2(new_n1189_), .ZN(new_n1358_));
  NAND3_X1  g1230(.A1(new_n1344_), .A2(new_n1351_), .A3(new_n1346_), .ZN(new_n1359_));
  NAND3_X1  g1231(.A1(new_n1357_), .A2(new_n1358_), .A3(new_n1359_), .ZN(new_n1360_));
  AOI21_X1  g1232(.A(new_n1226_), .B1(new_n1354_), .B2(new_n1360_), .ZN(new_n1361_));
  INV_X1    g1233(.A(new_n1361_), .ZN(new_n1362_));
  NAND3_X1  g1234(.A1(new_n1354_), .A2(new_n1360_), .A3(new_n1224_), .ZN(new_n1363_));
  NAND3_X1  g1235(.A1(new_n1223_), .A2(new_n1362_), .A3(new_n1363_), .ZN(new_n1364_));
  NAND3_X1  g1236(.A1(new_n1354_), .A2(new_n1360_), .A3(new_n1226_), .ZN(new_n1365_));
  INV_X1    g1237(.A(new_n1365_), .ZN(new_n1366_));
  OAI211_X1 g1238(.A(new_n1203_), .B(new_n1199_), .C1(new_n1361_), .C2(new_n1366_), .ZN(new_n1367_));
  NAND2_X1  g1239(.A1(G35gat), .A2(G494gat), .ZN(new_n1368_));
  NAND3_X1  g1240(.A1(new_n1364_), .A2(new_n1367_), .A3(new_n1368_), .ZN(new_n1369_));
  NAND2_X1  g1241(.A1(new_n1364_), .A2(new_n1367_), .ZN(new_n1370_));
  NAND3_X1  g1242(.A1(new_n1370_), .A2(G35gat), .A3(G494gat), .ZN(new_n1371_));
  AOI21_X1  g1243(.A(new_n1222_), .B1(new_n1369_), .B2(new_n1371_), .ZN(new_n1372_));
  INV_X1    g1244(.A(new_n1372_), .ZN(new_n1373_));
  NOR2_X1   g1245(.A1(new_n132_), .A2(new_n1218_), .ZN(new_n1374_));
  INV_X1    g1246(.A(new_n1374_), .ZN(new_n1375_));
  NAND3_X1  g1247(.A1(new_n1222_), .A2(new_n1371_), .A3(new_n1369_), .ZN(new_n1376_));
  NAND3_X1  g1248(.A1(new_n1373_), .A2(new_n1375_), .A3(new_n1376_), .ZN(new_n1377_));
  INV_X1    g1249(.A(new_n1376_), .ZN(new_n1378_));
  OAI21_X1  g1250(.A(new_n1374_), .B1(new_n1378_), .B2(new_n1372_), .ZN(new_n1379_));
  AOI21_X1  g1251(.A(new_n1221_), .B1(new_n1377_), .B2(new_n1379_), .ZN(new_n1380_));
  INV_X1    g1252(.A(new_n1380_), .ZN(new_n1381_));
  NAND3_X1  g1253(.A1(new_n1221_), .A2(new_n1377_), .A3(new_n1379_), .ZN(new_n1382_));
  NAND2_X1  g1254(.A1(new_n1381_), .A2(new_n1382_), .ZN(new_n1383_));
  INV_X1    g1255(.A(G528gat), .ZN(new_n1384_));
  NOR2_X1   g1256(.A1(new_n129_), .A2(new_n1384_), .ZN(new_n1385_));
  NAND2_X1  g1257(.A1(new_n1383_), .A2(new_n1385_), .ZN(new_n1386_));
  INV_X1    g1258(.A(new_n1385_), .ZN(new_n1387_));
  NAND3_X1  g1259(.A1(new_n1381_), .A2(new_n1387_), .A3(new_n1382_), .ZN(new_n1388_));
  NAND2_X1  g1260(.A1(new_n1386_), .A2(new_n1388_), .ZN(G6123gat));
  OAI21_X1  g1261(.A(new_n1376_), .B1(new_n1372_), .B2(new_n1374_), .ZN(new_n1390_));
  NAND3_X1  g1262(.A1(new_n1223_), .A2(new_n1362_), .A3(new_n1365_), .ZN(new_n1391_));
  AND2_X1   g1263(.A1(new_n1369_), .A2(new_n1391_), .ZN(new_n1392_));
  NOR2_X1   g1264(.A1(new_n165_), .A2(new_n1057_), .ZN(new_n1393_));
  NOR2_X1   g1265(.A1(new_n166_), .A2(new_n890_), .ZN(new_n1394_));
  NAND2_X1  g1266(.A1(new_n1359_), .A2(new_n1351_), .ZN(new_n1395_));
  AND3_X1   g1267(.A1(new_n1336_), .A2(new_n1339_), .A3(new_n1340_), .ZN(new_n1396_));
  AOI21_X1  g1268(.A(new_n1396_), .B1(new_n1335_), .B2(new_n1333_), .ZN(new_n1397_));
  AOI21_X1  g1269(.A(new_n1337_), .B1(new_n1321_), .B2(new_n1319_), .ZN(new_n1398_));
  NAND2_X1  g1270(.A1(new_n1309_), .A2(new_n1300_), .ZN(new_n1399_));
  NOR2_X1   g1271(.A1(new_n542_), .A2(new_n363_), .ZN(new_n1400_));
  INV_X1    g1272(.A(new_n1400_), .ZN(new_n1401_));
  NAND2_X1  g1273(.A1(new_n1267_), .A2(new_n1274_), .ZN(new_n1402_));
  NAND2_X1  g1274(.A1(new_n1402_), .A2(new_n1273_), .ZN(new_n1403_));
  AOI21_X1  g1275(.A(new_n1252_), .B1(new_n1245_), .B2(new_n1247_), .ZN(new_n1404_));
  AOI21_X1  g1276(.A(new_n1404_), .B1(new_n1259_), .B2(new_n1262_), .ZN(new_n1405_));
  INV_X1    g1277(.A(G222gat), .ZN(new_n1406_));
  NOR2_X1   g1278(.A1(new_n1406_), .A2(new_n159_), .ZN(new_n1407_));
  NAND3_X1  g1279(.A1(new_n1071_), .A2(G256gat), .A3(G290gat), .ZN(new_n1408_));
  NAND2_X1  g1280(.A1(G239gat), .A2(G307gat), .ZN(new_n1409_));
  XNOR2_X1  g1281(.A(new_n1408_), .B(new_n1409_), .ZN(new_n1410_));
  NOR2_X1   g1282(.A1(new_n1240_), .A2(new_n1254_), .ZN(new_n1411_));
  INV_X1    g1283(.A(new_n1411_), .ZN(new_n1412_));
  NAND3_X1  g1284(.A1(new_n1256_), .A2(new_n1410_), .A3(new_n1412_), .ZN(new_n1413_));
  AOI21_X1  g1285(.A(new_n1411_), .B1(new_n1242_), .B2(new_n1243_), .ZN(new_n1414_));
  OAI211_X1 g1286(.A(new_n1407_), .B(new_n1413_), .C1(new_n1414_), .C2(new_n1410_), .ZN(new_n1415_));
  INV_X1    g1287(.A(new_n1407_), .ZN(new_n1416_));
  INV_X1    g1288(.A(new_n1410_), .ZN(new_n1417_));
  NAND3_X1  g1289(.A1(new_n1256_), .A2(new_n1417_), .A3(new_n1412_), .ZN(new_n1418_));
  OAI211_X1 g1290(.A(new_n1416_), .B(new_n1418_), .C1(new_n1414_), .C2(new_n1417_), .ZN(new_n1419_));
  NAND2_X1  g1291(.A1(new_n1415_), .A2(new_n1419_), .ZN(new_n1420_));
  NAND2_X1  g1292(.A1(new_n1405_), .A2(new_n1420_), .ZN(new_n1421_));
  NOR2_X1   g1293(.A1(new_n1260_), .A2(new_n198_), .ZN(new_n1422_));
  INV_X1    g1294(.A(new_n1422_), .ZN(new_n1423_));
  OAI211_X1 g1295(.A(new_n1415_), .B(new_n1419_), .C1(new_n1272_), .C2(new_n1404_), .ZN(new_n1424_));
  NAND3_X1  g1296(.A1(new_n1421_), .A2(new_n1423_), .A3(new_n1424_), .ZN(new_n1425_));
  INV_X1    g1297(.A(new_n1425_), .ZN(new_n1426_));
  AOI21_X1  g1298(.A(new_n1423_), .B1(new_n1421_), .B2(new_n1424_), .ZN(new_n1427_));
  OAI21_X1  g1299(.A(new_n1403_), .B1(new_n1426_), .B2(new_n1427_), .ZN(new_n1428_));
  INV_X1    g1300(.A(new_n1427_), .ZN(new_n1429_));
  AOI21_X1  g1301(.A(new_n1269_), .B1(new_n1274_), .B2(new_n1267_), .ZN(new_n1430_));
  NAND3_X1  g1302(.A1(new_n1429_), .A2(new_n1425_), .A3(new_n1430_), .ZN(new_n1431_));
  NOR2_X1   g1303(.A1(new_n1084_), .A2(new_n276_), .ZN(new_n1432_));
  INV_X1    g1304(.A(new_n1432_), .ZN(new_n1433_));
  AND3_X1   g1305(.A1(new_n1428_), .A2(new_n1431_), .A3(new_n1433_), .ZN(new_n1434_));
  AOI21_X1  g1306(.A(new_n1433_), .B1(new_n1428_), .B2(new_n1431_), .ZN(new_n1435_));
  OR2_X1    g1307(.A1(new_n1434_), .A2(new_n1435_), .ZN(new_n1436_));
  NOR2_X1   g1308(.A1(new_n1107_), .A2(new_n1276_), .ZN(new_n1437_));
  NAND2_X1  g1309(.A1(new_n1280_), .A2(new_n1281_), .ZN(new_n1438_));
  NOR2_X1   g1310(.A1(new_n1437_), .A2(new_n1438_), .ZN(new_n1439_));
  INV_X1    g1311(.A(new_n1439_), .ZN(new_n1440_));
  NAND3_X1  g1312(.A1(new_n1290_), .A2(new_n1436_), .A3(new_n1440_), .ZN(new_n1441_));
  NOR2_X1   g1313(.A1(new_n1434_), .A2(new_n1435_), .ZN(new_n1442_));
  OAI21_X1  g1314(.A(new_n1442_), .B1(new_n1286_), .B2(new_n1439_), .ZN(new_n1443_));
  NOR2_X1   g1315(.A1(new_n543_), .A2(new_n289_), .ZN(new_n1444_));
  INV_X1    g1316(.A(new_n1444_), .ZN(new_n1445_));
  AND3_X1   g1317(.A1(new_n1441_), .A2(new_n1443_), .A3(new_n1445_), .ZN(new_n1446_));
  AOI21_X1  g1318(.A(new_n1445_), .B1(new_n1441_), .B2(new_n1443_), .ZN(new_n1447_));
  NOR2_X1   g1319(.A1(new_n1446_), .A2(new_n1447_), .ZN(new_n1448_));
  NAND2_X1  g1320(.A1(new_n1297_), .A2(new_n1292_), .ZN(new_n1449_));
  NAND2_X1  g1321(.A1(new_n1448_), .A2(new_n1449_), .ZN(new_n1450_));
  OAI211_X1 g1322(.A(new_n1297_), .B(new_n1292_), .C1(new_n1446_), .C2(new_n1447_), .ZN(new_n1451_));
  AOI21_X1  g1323(.A(new_n1401_), .B1(new_n1450_), .B2(new_n1451_), .ZN(new_n1452_));
  INV_X1    g1324(.A(new_n1452_), .ZN(new_n1453_));
  NAND3_X1  g1325(.A1(new_n1450_), .A2(new_n1401_), .A3(new_n1451_), .ZN(new_n1454_));
  NAND3_X1  g1326(.A1(new_n1399_), .A2(new_n1453_), .A3(new_n1454_), .ZN(new_n1455_));
  AND3_X1   g1327(.A1(new_n1450_), .A2(new_n1401_), .A3(new_n1451_), .ZN(new_n1456_));
  OAI211_X1 g1328(.A(new_n1300_), .B(new_n1309_), .C1(new_n1456_), .C2(new_n1452_), .ZN(new_n1457_));
  NOR2_X1   g1329(.A1(new_n377_), .A2(new_n443_), .ZN(new_n1458_));
  INV_X1    g1330(.A(new_n1458_), .ZN(new_n1459_));
  AND3_X1   g1331(.A1(new_n1455_), .A2(new_n1457_), .A3(new_n1459_), .ZN(new_n1460_));
  AOI21_X1  g1332(.A(new_n1459_), .B1(new_n1455_), .B2(new_n1457_), .ZN(new_n1461_));
  NOR2_X1   g1333(.A1(new_n1460_), .A2(new_n1461_), .ZN(new_n1462_));
  NAND2_X1  g1334(.A1(new_n1324_), .A2(new_n1311_), .ZN(new_n1463_));
  NAND2_X1  g1335(.A1(new_n1329_), .A2(new_n1463_), .ZN(new_n1464_));
  NAND2_X1  g1336(.A1(new_n1462_), .A2(new_n1464_), .ZN(new_n1465_));
  NOR2_X1   g1337(.A1(new_n300_), .A2(new_n533_), .ZN(new_n1466_));
  INV_X1    g1338(.A(new_n1466_), .ZN(new_n1467_));
  OAI211_X1 g1339(.A(new_n1329_), .B(new_n1463_), .C1(new_n1460_), .C2(new_n1461_), .ZN(new_n1468_));
  AND3_X1   g1340(.A1(new_n1465_), .A2(new_n1467_), .A3(new_n1468_), .ZN(new_n1469_));
  AOI21_X1  g1341(.A(new_n1467_), .B1(new_n1465_), .B2(new_n1468_), .ZN(new_n1470_));
  OAI21_X1  g1342(.A(new_n1398_), .B1(new_n1469_), .B2(new_n1470_), .ZN(new_n1471_));
  NAND2_X1  g1343(.A1(new_n1465_), .A2(new_n1468_), .ZN(new_n1472_));
  NAND2_X1  g1344(.A1(new_n1472_), .A2(new_n1466_), .ZN(new_n1473_));
  OAI21_X1  g1345(.A(new_n1330_), .B1(new_n1338_), .B2(new_n1320_), .ZN(new_n1474_));
  NAND3_X1  g1346(.A1(new_n1465_), .A2(new_n1467_), .A3(new_n1468_), .ZN(new_n1475_));
  NAND3_X1  g1347(.A1(new_n1473_), .A2(new_n1474_), .A3(new_n1475_), .ZN(new_n1476_));
  NOR2_X1   g1348(.A1(new_n243_), .A2(new_n648_), .ZN(new_n1477_));
  INV_X1    g1349(.A(new_n1477_), .ZN(new_n1478_));
  AND3_X1   g1350(.A1(new_n1471_), .A2(new_n1476_), .A3(new_n1478_), .ZN(new_n1479_));
  AOI21_X1  g1351(.A(new_n1478_), .B1(new_n1471_), .B2(new_n1476_), .ZN(new_n1480_));
  OAI21_X1  g1352(.A(new_n1397_), .B1(new_n1479_), .B2(new_n1480_), .ZN(new_n1481_));
  NOR3_X1   g1353(.A1(new_n1398_), .A2(new_n1469_), .A3(new_n1470_), .ZN(new_n1482_));
  AOI21_X1  g1354(.A(new_n1474_), .B1(new_n1473_), .B2(new_n1475_), .ZN(new_n1483_));
  OAI21_X1  g1355(.A(new_n1477_), .B1(new_n1482_), .B2(new_n1483_), .ZN(new_n1484_));
  AOI21_X1  g1356(.A(new_n1336_), .B1(new_n1340_), .B2(new_n1339_), .ZN(new_n1485_));
  OAI21_X1  g1357(.A(new_n1341_), .B1(new_n1485_), .B2(new_n1334_), .ZN(new_n1486_));
  NAND3_X1  g1358(.A1(new_n1471_), .A2(new_n1476_), .A3(new_n1478_), .ZN(new_n1487_));
  NAND3_X1  g1359(.A1(new_n1484_), .A2(new_n1486_), .A3(new_n1487_), .ZN(new_n1488_));
  NOR2_X1   g1360(.A1(new_n242_), .A2(new_n654_), .ZN(new_n1489_));
  INV_X1    g1361(.A(new_n1489_), .ZN(new_n1490_));
  AND3_X1   g1362(.A1(new_n1481_), .A2(new_n1488_), .A3(new_n1490_), .ZN(new_n1491_));
  AOI21_X1  g1363(.A(new_n1490_), .B1(new_n1481_), .B2(new_n1488_), .ZN(new_n1492_));
  NOR2_X1   g1364(.A1(new_n1491_), .A2(new_n1492_), .ZN(new_n1493_));
  NAND2_X1  g1365(.A1(new_n1359_), .A2(KEYINPUT41), .ZN(new_n1494_));
  AOI21_X1  g1366(.A(new_n1395_), .B1(new_n1493_), .B2(new_n1494_), .ZN(new_n1495_));
  NAND3_X1  g1367(.A1(new_n1481_), .A2(new_n1488_), .A3(new_n1490_), .ZN(new_n1496_));
  NAND2_X1  g1368(.A1(new_n1481_), .A2(new_n1488_), .ZN(new_n1497_));
  NAND2_X1  g1369(.A1(new_n1497_), .A2(new_n1489_), .ZN(new_n1498_));
  AND4_X1   g1370(.A1(new_n1395_), .A2(new_n1494_), .A3(new_n1496_), .A4(new_n1498_), .ZN(new_n1499_));
  OAI21_X1  g1371(.A(new_n1394_), .B1(new_n1495_), .B2(new_n1499_), .ZN(new_n1500_));
  NAND3_X1  g1372(.A1(new_n1494_), .A2(new_n1498_), .A3(new_n1496_), .ZN(new_n1501_));
  INV_X1    g1373(.A(new_n1395_), .ZN(new_n1502_));
  NAND2_X1  g1374(.A1(new_n1501_), .A2(new_n1502_), .ZN(new_n1503_));
  NAND3_X1  g1375(.A1(new_n1493_), .A2(new_n1395_), .A3(new_n1494_), .ZN(new_n1504_));
  INV_X1    g1376(.A(new_n1394_), .ZN(new_n1505_));
  NAND3_X1  g1377(.A1(new_n1503_), .A2(new_n1504_), .A3(new_n1505_), .ZN(new_n1506_));
  INV_X1    g1378(.A(KEYINPUT40), .ZN(new_n1507_));
  XNOR2_X1  g1379(.A(new_n1360_), .B(new_n1507_), .ZN(new_n1508_));
  NAND4_X1  g1380(.A1(new_n1500_), .A2(new_n1365_), .A3(new_n1506_), .A4(new_n1508_), .ZN(new_n1509_));
  NOR3_X1   g1381(.A1(new_n1495_), .A2(new_n1499_), .A3(new_n1394_), .ZN(new_n1510_));
  AOI21_X1  g1382(.A(new_n1505_), .B1(new_n1503_), .B2(new_n1504_), .ZN(new_n1511_));
  NOR2_X1   g1383(.A1(new_n1510_), .A2(new_n1511_), .ZN(new_n1512_));
  XNOR2_X1  g1384(.A(new_n1360_), .B(KEYINPUT40), .ZN(new_n1513_));
  NAND2_X1  g1385(.A1(new_n1363_), .A2(KEYINPUT42), .ZN(new_n1514_));
  INV_X1    g1386(.A(KEYINPUT42), .ZN(new_n1515_));
  NAND4_X1  g1387(.A1(new_n1354_), .A2(new_n1360_), .A3(new_n1515_), .A4(new_n1224_), .ZN(new_n1516_));
  AOI21_X1  g1388(.A(new_n1513_), .B1(new_n1514_), .B2(new_n1516_), .ZN(new_n1517_));
  OAI211_X1 g1389(.A(new_n1393_), .B(new_n1509_), .C1(new_n1512_), .C2(new_n1517_), .ZN(new_n1518_));
  INV_X1    g1390(.A(new_n1518_), .ZN(new_n1519_));
  NAND2_X1  g1391(.A1(new_n1514_), .A2(new_n1516_), .ZN(new_n1520_));
  NAND2_X1  g1392(.A1(new_n1520_), .A2(new_n1508_), .ZN(new_n1521_));
  NAND2_X1  g1393(.A1(new_n1500_), .A2(new_n1506_), .ZN(new_n1522_));
  NAND2_X1  g1394(.A1(new_n1521_), .A2(new_n1522_), .ZN(new_n1523_));
  AOI21_X1  g1395(.A(new_n1393_), .B1(new_n1523_), .B2(new_n1509_), .ZN(new_n1524_));
  OAI21_X1  g1396(.A(new_n1392_), .B1(new_n1519_), .B2(new_n1524_), .ZN(new_n1525_));
  INV_X1    g1397(.A(new_n1393_), .ZN(new_n1526_));
  AOI22_X1  g1398(.A1(new_n1520_), .A2(new_n1508_), .B1(new_n1500_), .B2(new_n1506_), .ZN(new_n1527_));
  NOR2_X1   g1399(.A1(new_n1352_), .A2(new_n1353_), .ZN(new_n1528_));
  AOI21_X1  g1400(.A(KEYINPUT40), .B1(new_n1528_), .B2(new_n1358_), .ZN(new_n1529_));
  NOR2_X1   g1401(.A1(new_n1360_), .A2(new_n1507_), .ZN(new_n1530_));
  OAI21_X1  g1402(.A(new_n1365_), .B1(new_n1529_), .B2(new_n1530_), .ZN(new_n1531_));
  NOR3_X1   g1403(.A1(new_n1510_), .A2(new_n1531_), .A3(new_n1511_), .ZN(new_n1532_));
  OAI21_X1  g1404(.A(new_n1526_), .B1(new_n1527_), .B2(new_n1532_), .ZN(new_n1533_));
  NAND2_X1  g1405(.A1(new_n1369_), .A2(new_n1391_), .ZN(new_n1534_));
  NAND3_X1  g1406(.A1(new_n1533_), .A2(new_n1534_), .A3(new_n1518_), .ZN(new_n1535_));
  NAND2_X1  g1407(.A1(new_n1525_), .A2(new_n1535_), .ZN(new_n1536_));
  NOR2_X1   g1408(.A1(new_n218_), .A2(new_n1218_), .ZN(new_n1537_));
  NAND2_X1  g1409(.A1(new_n1536_), .A2(new_n1537_), .ZN(new_n1538_));
  OAI211_X1 g1410(.A(new_n1525_), .B(new_n1535_), .C1(new_n218_), .C2(new_n1218_), .ZN(new_n1539_));
  AOI21_X1  g1411(.A(new_n1390_), .B1(new_n1538_), .B2(new_n1539_), .ZN(new_n1540_));
  INV_X1    g1412(.A(new_n1540_), .ZN(new_n1541_));
  NOR2_X1   g1413(.A1(new_n132_), .A2(new_n1384_), .ZN(new_n1542_));
  INV_X1    g1414(.A(new_n1542_), .ZN(new_n1543_));
  AND3_X1   g1415(.A1(new_n1538_), .A2(new_n1390_), .A3(new_n1539_), .ZN(new_n1544_));
  INV_X1    g1416(.A(new_n1544_), .ZN(new_n1545_));
  NAND3_X1  g1417(.A1(new_n1541_), .A2(new_n1543_), .A3(new_n1545_), .ZN(new_n1546_));
  OAI21_X1  g1418(.A(new_n1542_), .B1(new_n1544_), .B2(new_n1540_), .ZN(new_n1547_));
  NAND2_X1  g1419(.A1(new_n1546_), .A2(new_n1547_), .ZN(new_n1548_));
  OAI21_X1  g1420(.A(new_n1382_), .B1(new_n1380_), .B2(new_n1385_), .ZN(new_n1549_));
  XNOR2_X1  g1421(.A(new_n1548_), .B(new_n1549_), .ZN(G6150gat));
  AOI21_X1  g1422(.A(new_n1544_), .B1(new_n1541_), .B2(new_n1543_), .ZN(new_n1551_));
  NOR3_X1   g1423(.A1(new_n1397_), .A2(new_n1479_), .A3(new_n1480_), .ZN(new_n1552_));
  AOI21_X1  g1424(.A(new_n1552_), .B1(new_n1490_), .B2(new_n1481_), .ZN(new_n1553_));
  AOI21_X1  g1425(.A(new_n1482_), .B1(new_n1478_), .B2(new_n1471_), .ZN(new_n1554_));
  INV_X1    g1426(.A(KEYINPUT45), .ZN(new_n1555_));
  NAND2_X1  g1427(.A1(new_n1464_), .A2(new_n1555_), .ZN(new_n1556_));
  INV_X1    g1428(.A(KEYINPUT44), .ZN(new_n1557_));
  OAI21_X1  g1429(.A(new_n1557_), .B1(new_n1460_), .B2(new_n1461_), .ZN(new_n1558_));
  INV_X1    g1430(.A(new_n1461_), .ZN(new_n1559_));
  NAND3_X1  g1431(.A1(new_n1455_), .A2(new_n1457_), .A3(new_n1459_), .ZN(new_n1560_));
  NAND3_X1  g1432(.A1(new_n1559_), .A2(KEYINPUT44), .A3(new_n1560_), .ZN(new_n1561_));
  NAND3_X1  g1433(.A1(new_n1329_), .A2(KEYINPUT45), .A3(new_n1463_), .ZN(new_n1562_));
  NAND4_X1  g1434(.A1(new_n1556_), .A2(new_n1558_), .A3(new_n1561_), .A4(new_n1562_), .ZN(new_n1563_));
  NOR2_X1   g1435(.A1(new_n377_), .A2(new_n533_), .ZN(new_n1564_));
  AND3_X1   g1436(.A1(new_n1399_), .A2(new_n1453_), .A3(new_n1454_), .ZN(new_n1565_));
  AOI21_X1  g1437(.A(new_n1565_), .B1(new_n1459_), .B2(new_n1457_), .ZN(new_n1566_));
  NOR2_X1   g1438(.A1(new_n1084_), .A2(new_n289_), .ZN(new_n1567_));
  NOR3_X1   g1439(.A1(new_n1426_), .A2(new_n1403_), .A3(new_n1427_), .ZN(new_n1568_));
  AOI21_X1  g1440(.A(new_n1568_), .B1(new_n1433_), .B2(new_n1428_), .ZN(new_n1569_));
  NAND2_X1  g1441(.A1(new_n1425_), .A2(new_n1424_), .ZN(new_n1570_));
  NOR2_X1   g1442(.A1(new_n1406_), .A2(new_n198_), .ZN(new_n1571_));
  INV_X1    g1443(.A(new_n1571_), .ZN(new_n1572_));
  NAND2_X1  g1444(.A1(new_n1418_), .A2(new_n1416_), .ZN(new_n1573_));
  NAND4_X1  g1445(.A1(new_n1071_), .A2(new_n1409_), .A3(G256gat), .A4(G290gat), .ZN(new_n1574_));
  NAND2_X1  g1446(.A1(new_n1574_), .A2(G290gat), .ZN(new_n1575_));
  AOI21_X1  g1447(.A(new_n1232_), .B1(new_n1575_), .B2(new_n150_), .ZN(new_n1576_));
  OAI21_X1  g1448(.A(new_n1576_), .B1(new_n133_), .B2(new_n1409_), .ZN(new_n1577_));
  INV_X1    g1449(.A(G239gat), .ZN(new_n1578_));
  NOR2_X1   g1450(.A1(new_n1578_), .A2(new_n159_), .ZN(new_n1579_));
  NAND2_X1  g1451(.A1(new_n1577_), .A2(new_n1579_), .ZN(new_n1580_));
  OAI221_X1 g1452(.A(new_n1576_), .B1(new_n1578_), .B2(new_n159_), .C1(new_n133_), .C2(new_n1409_), .ZN(new_n1581_));
  NAND2_X1  g1453(.A1(new_n1580_), .A2(new_n1581_), .ZN(new_n1582_));
  OAI211_X1 g1454(.A(new_n1573_), .B(new_n1582_), .C1(new_n1417_), .C2(new_n1414_), .ZN(new_n1583_));
  NOR2_X1   g1455(.A1(new_n1414_), .A2(new_n1417_), .ZN(new_n1584_));
  OAI21_X1  g1456(.A(new_n1413_), .B1(new_n1414_), .B2(new_n1410_), .ZN(new_n1585_));
  AOI21_X1  g1457(.A(new_n1584_), .B1(new_n1585_), .B2(new_n1416_), .ZN(new_n1586_));
  OAI211_X1 g1458(.A(new_n1572_), .B(new_n1583_), .C1(new_n1586_), .C2(new_n1582_), .ZN(new_n1587_));
  INV_X1    g1459(.A(new_n1582_), .ZN(new_n1588_));
  OAI211_X1 g1460(.A(new_n1588_), .B(new_n1573_), .C1(new_n1417_), .C2(new_n1414_), .ZN(new_n1589_));
  OAI211_X1 g1461(.A(new_n1589_), .B(new_n1571_), .C1(new_n1586_), .C2(new_n1588_), .ZN(new_n1590_));
  AND2_X1   g1462(.A1(new_n1587_), .A2(new_n1590_), .ZN(new_n1591_));
  NAND2_X1  g1463(.A1(new_n1570_), .A2(new_n1591_), .ZN(new_n1592_));
  NAND2_X1  g1464(.A1(new_n1587_), .A2(new_n1590_), .ZN(new_n1593_));
  NAND3_X1  g1465(.A1(new_n1593_), .A2(new_n1425_), .A3(new_n1424_), .ZN(new_n1594_));
  NOR2_X1   g1466(.A1(new_n1260_), .A2(new_n276_), .ZN(new_n1595_));
  INV_X1    g1467(.A(new_n1595_), .ZN(new_n1596_));
  AND3_X1   g1468(.A1(new_n1592_), .A2(new_n1594_), .A3(new_n1596_), .ZN(new_n1597_));
  AOI21_X1  g1469(.A(new_n1596_), .B1(new_n1592_), .B2(new_n1594_), .ZN(new_n1598_));
  NOR3_X1   g1470(.A1(new_n1569_), .A2(new_n1597_), .A3(new_n1598_), .ZN(new_n1599_));
  AOI21_X1  g1471(.A(new_n1430_), .B1(new_n1429_), .B2(new_n1425_), .ZN(new_n1600_));
  OAI21_X1  g1472(.A(new_n1431_), .B1(new_n1600_), .B2(new_n1432_), .ZN(new_n1601_));
  INV_X1    g1473(.A(new_n1598_), .ZN(new_n1602_));
  NAND3_X1  g1474(.A1(new_n1592_), .A2(new_n1594_), .A3(new_n1596_), .ZN(new_n1603_));
  AOI21_X1  g1475(.A(new_n1601_), .B1(new_n1602_), .B2(new_n1603_), .ZN(new_n1604_));
  OAI21_X1  g1476(.A(new_n1567_), .B1(new_n1599_), .B2(new_n1604_), .ZN(new_n1605_));
  OAI21_X1  g1477(.A(new_n1569_), .B1(new_n1597_), .B2(new_n1598_), .ZN(new_n1606_));
  NAND3_X1  g1478(.A1(new_n1602_), .A2(new_n1601_), .A3(new_n1603_), .ZN(new_n1607_));
  INV_X1    g1479(.A(new_n1567_), .ZN(new_n1608_));
  NAND3_X1  g1480(.A1(new_n1606_), .A2(new_n1607_), .A3(new_n1608_), .ZN(new_n1609_));
  AND2_X1   g1481(.A1(new_n1605_), .A2(new_n1609_), .ZN(new_n1610_));
  NOR3_X1   g1482(.A1(new_n1286_), .A2(new_n1442_), .A3(new_n1439_), .ZN(new_n1611_));
  OAI21_X1  g1483(.A(new_n1443_), .B1(new_n1611_), .B2(new_n1444_), .ZN(new_n1612_));
  NAND2_X1  g1484(.A1(new_n1610_), .A2(new_n1612_), .ZN(new_n1613_));
  NAND3_X1  g1485(.A1(new_n1441_), .A2(new_n1443_), .A3(new_n1445_), .ZN(new_n1614_));
  NAND2_X1  g1486(.A1(new_n1605_), .A2(new_n1609_), .ZN(new_n1615_));
  NAND3_X1  g1487(.A1(new_n1614_), .A2(new_n1615_), .A3(new_n1443_), .ZN(new_n1616_));
  NOR2_X1   g1488(.A1(new_n543_), .A2(new_n363_), .ZN(new_n1617_));
  INV_X1    g1489(.A(new_n1617_), .ZN(new_n1618_));
  AND3_X1   g1490(.A1(new_n1613_), .A2(new_n1616_), .A3(new_n1618_), .ZN(new_n1619_));
  AOI21_X1  g1491(.A(new_n1618_), .B1(new_n1613_), .B2(new_n1616_), .ZN(new_n1620_));
  OAI211_X1 g1492(.A(new_n1454_), .B(new_n1450_), .C1(new_n1619_), .C2(new_n1620_), .ZN(new_n1621_));
  INV_X1    g1493(.A(new_n1451_), .ZN(new_n1622_));
  OAI21_X1  g1494(.A(new_n1450_), .B1(new_n1622_), .B2(new_n1400_), .ZN(new_n1623_));
  NOR2_X1   g1495(.A1(new_n1619_), .A2(new_n1620_), .ZN(new_n1624_));
  NAND2_X1  g1496(.A1(new_n1623_), .A2(new_n1624_), .ZN(new_n1625_));
  NAND2_X1  g1497(.A1(new_n1621_), .A2(new_n1625_), .ZN(new_n1626_));
  NOR2_X1   g1498(.A1(new_n542_), .A2(new_n443_), .ZN(new_n1627_));
  NAND2_X1  g1499(.A1(new_n1626_), .A2(new_n1627_), .ZN(new_n1628_));
  INV_X1    g1500(.A(new_n1627_), .ZN(new_n1629_));
  NAND3_X1  g1501(.A1(new_n1621_), .A2(new_n1625_), .A3(new_n1629_), .ZN(new_n1630_));
  NAND2_X1  g1502(.A1(new_n1628_), .A2(new_n1630_), .ZN(new_n1631_));
  NOR2_X1   g1503(.A1(new_n1566_), .A2(new_n1631_), .ZN(new_n1632_));
  AND3_X1   g1504(.A1(new_n1621_), .A2(new_n1625_), .A3(new_n1629_), .ZN(new_n1633_));
  AOI21_X1  g1505(.A(new_n1629_), .B1(new_n1621_), .B2(new_n1625_), .ZN(new_n1634_));
  NOR2_X1   g1506(.A1(new_n1633_), .A2(new_n1634_), .ZN(new_n1635_));
  INV_X1    g1507(.A(new_n1457_), .ZN(new_n1636_));
  OAI21_X1  g1508(.A(new_n1455_), .B1(new_n1636_), .B2(new_n1458_), .ZN(new_n1637_));
  NOR2_X1   g1509(.A1(new_n1635_), .A2(new_n1637_), .ZN(new_n1638_));
  OAI21_X1  g1510(.A(new_n1564_), .B1(new_n1632_), .B2(new_n1638_), .ZN(new_n1639_));
  NAND2_X1  g1511(.A1(new_n1566_), .A2(new_n1631_), .ZN(new_n1640_));
  NAND2_X1  g1512(.A1(new_n1635_), .A2(new_n1637_), .ZN(new_n1641_));
  INV_X1    g1513(.A(new_n1564_), .ZN(new_n1642_));
  NAND3_X1  g1514(.A1(new_n1640_), .A2(new_n1641_), .A3(new_n1642_), .ZN(new_n1643_));
  NAND2_X1  g1515(.A1(new_n1639_), .A2(new_n1643_), .ZN(new_n1644_));
  OAI211_X1 g1516(.A(new_n1475_), .B(new_n1563_), .C1(new_n1644_), .C2(KEYINPUT43), .ZN(new_n1645_));
  NAND2_X1  g1517(.A1(new_n1563_), .A2(new_n1475_), .ZN(new_n1646_));
  NAND2_X1  g1518(.A1(new_n1563_), .A2(KEYINPUT43), .ZN(new_n1647_));
  AND3_X1   g1519(.A1(new_n1640_), .A2(new_n1641_), .A3(new_n1642_), .ZN(new_n1648_));
  AOI21_X1  g1520(.A(new_n1642_), .B1(new_n1640_), .B2(new_n1641_), .ZN(new_n1649_));
  NOR2_X1   g1521(.A1(new_n1648_), .A2(new_n1649_), .ZN(new_n1650_));
  NAND3_X1  g1522(.A1(new_n1646_), .A2(new_n1647_), .A3(new_n1650_), .ZN(new_n1651_));
  NOR2_X1   g1523(.A1(new_n300_), .A2(new_n648_), .ZN(new_n1652_));
  INV_X1    g1524(.A(new_n1652_), .ZN(new_n1653_));
  AND3_X1   g1525(.A1(new_n1645_), .A2(new_n1651_), .A3(new_n1653_), .ZN(new_n1654_));
  AOI21_X1  g1526(.A(new_n1653_), .B1(new_n1645_), .B2(new_n1651_), .ZN(new_n1655_));
  OAI21_X1  g1527(.A(new_n1554_), .B1(new_n1654_), .B2(new_n1655_), .ZN(new_n1656_));
  NAND2_X1  g1528(.A1(new_n1645_), .A2(new_n1651_), .ZN(new_n1657_));
  NAND2_X1  g1529(.A1(new_n1657_), .A2(new_n1652_), .ZN(new_n1658_));
  NAND2_X1  g1530(.A1(new_n1487_), .A2(new_n1476_), .ZN(new_n1659_));
  NAND3_X1  g1531(.A1(new_n1645_), .A2(new_n1651_), .A3(new_n1653_), .ZN(new_n1660_));
  NAND3_X1  g1532(.A1(new_n1658_), .A2(new_n1659_), .A3(new_n1660_), .ZN(new_n1661_));
  NOR2_X1   g1533(.A1(new_n243_), .A2(new_n654_), .ZN(new_n1662_));
  INV_X1    g1534(.A(new_n1662_), .ZN(new_n1663_));
  AND3_X1   g1535(.A1(new_n1656_), .A2(new_n1661_), .A3(new_n1663_), .ZN(new_n1664_));
  AOI21_X1  g1536(.A(new_n1663_), .B1(new_n1656_), .B2(new_n1661_), .ZN(new_n1665_));
  OAI21_X1  g1537(.A(new_n1553_), .B1(new_n1664_), .B2(new_n1665_), .ZN(new_n1666_));
  NOR3_X1   g1538(.A1(new_n1654_), .A2(new_n1554_), .A3(new_n1655_), .ZN(new_n1667_));
  AOI21_X1  g1539(.A(new_n1659_), .B1(new_n1658_), .B2(new_n1660_), .ZN(new_n1668_));
  OAI21_X1  g1540(.A(new_n1662_), .B1(new_n1667_), .B2(new_n1668_), .ZN(new_n1669_));
  NAND2_X1  g1541(.A1(new_n1496_), .A2(new_n1488_), .ZN(new_n1670_));
  NAND3_X1  g1542(.A1(new_n1656_), .A2(new_n1661_), .A3(new_n1663_), .ZN(new_n1671_));
  NAND3_X1  g1543(.A1(new_n1669_), .A2(new_n1670_), .A3(new_n1671_), .ZN(new_n1672_));
  NAND2_X1  g1544(.A1(G86gat), .A2(G477gat), .ZN(new_n1673_));
  XNOR2_X1  g1545(.A(new_n1673_), .B(KEYINPUT46), .ZN(new_n1674_));
  AND3_X1   g1546(.A1(new_n1666_), .A2(new_n1672_), .A3(new_n1674_), .ZN(new_n1675_));
  AOI21_X1  g1547(.A(new_n1674_), .B1(new_n1666_), .B2(new_n1672_), .ZN(new_n1676_));
  NOR2_X1   g1548(.A1(new_n1675_), .A2(new_n1676_), .ZN(new_n1677_));
  NAND2_X1  g1549(.A1(new_n1493_), .A2(new_n1395_), .ZN(new_n1678_));
  NAND2_X1  g1550(.A1(new_n1506_), .A2(new_n1678_), .ZN(new_n1679_));
  NAND2_X1  g1551(.A1(new_n1677_), .A2(new_n1679_), .ZN(new_n1680_));
  NOR2_X1   g1552(.A1(new_n166_), .A2(new_n1057_), .ZN(new_n1681_));
  INV_X1    g1553(.A(new_n1681_), .ZN(new_n1682_));
  OAI211_X1 g1554(.A(new_n1506_), .B(new_n1678_), .C1(new_n1675_), .C2(new_n1676_), .ZN(new_n1683_));
  NAND3_X1  g1555(.A1(new_n1680_), .A2(new_n1682_), .A3(new_n1683_), .ZN(new_n1684_));
  NAND2_X1  g1556(.A1(new_n1680_), .A2(new_n1683_), .ZN(new_n1685_));
  NAND2_X1  g1557(.A1(new_n1685_), .A2(new_n1681_), .ZN(new_n1686_));
  NOR2_X1   g1558(.A1(new_n1517_), .A2(new_n1522_), .ZN(new_n1687_));
  OAI211_X1 g1559(.A(new_n1684_), .B(new_n1686_), .C1(new_n1524_), .C2(new_n1687_), .ZN(new_n1688_));
  NOR2_X1   g1560(.A1(new_n165_), .A2(new_n1218_), .ZN(new_n1689_));
  INV_X1    g1561(.A(new_n1687_), .ZN(new_n1690_));
  AND3_X1   g1562(.A1(new_n1680_), .A2(new_n1682_), .A3(new_n1683_), .ZN(new_n1691_));
  AOI21_X1  g1563(.A(new_n1682_), .B1(new_n1680_), .B2(new_n1683_), .ZN(new_n1692_));
  OAI211_X1 g1564(.A(new_n1533_), .B(new_n1690_), .C1(new_n1691_), .C2(new_n1692_), .ZN(new_n1693_));
  NAND3_X1  g1565(.A1(new_n1688_), .A2(new_n1689_), .A3(new_n1693_), .ZN(new_n1694_));
  INV_X1    g1566(.A(KEYINPUT47), .ZN(new_n1695_));
  NAND2_X1  g1567(.A1(new_n1694_), .A2(new_n1695_), .ZN(new_n1696_));
  NAND2_X1  g1568(.A1(new_n1688_), .A2(new_n1693_), .ZN(new_n1697_));
  INV_X1    g1569(.A(new_n1689_), .ZN(new_n1698_));
  NAND2_X1  g1570(.A1(new_n1697_), .A2(new_n1698_), .ZN(new_n1699_));
  NAND4_X1  g1571(.A1(new_n1688_), .A2(new_n1693_), .A3(KEYINPUT47), .A4(new_n1689_), .ZN(new_n1700_));
  NAND3_X1  g1572(.A1(new_n1696_), .A2(new_n1699_), .A3(new_n1700_), .ZN(new_n1701_));
  AOI21_X1  g1573(.A(new_n1534_), .B1(new_n1533_), .B2(new_n1518_), .ZN(new_n1702_));
  OAI21_X1  g1574(.A(new_n1535_), .B1(new_n1702_), .B2(new_n1537_), .ZN(new_n1703_));
  INV_X1    g1575(.A(new_n1703_), .ZN(new_n1704_));
  NAND2_X1  g1576(.A1(new_n1701_), .A2(new_n1704_), .ZN(new_n1705_));
  NOR2_X1   g1577(.A1(new_n218_), .A2(new_n1384_), .ZN(new_n1706_));
  AND2_X1   g1578(.A1(new_n1703_), .A2(new_n1694_), .ZN(new_n1707_));
  NAND2_X1  g1579(.A1(new_n1707_), .A2(new_n1699_), .ZN(new_n1708_));
  AND3_X1   g1580(.A1(new_n1705_), .A2(new_n1706_), .A3(new_n1708_), .ZN(new_n1709_));
  AOI21_X1  g1581(.A(new_n1706_), .B1(new_n1705_), .B2(new_n1708_), .ZN(new_n1710_));
  OAI21_X1  g1582(.A(new_n1551_), .B1(new_n1709_), .B2(new_n1710_), .ZN(new_n1711_));
  NAND2_X1  g1583(.A1(new_n1705_), .A2(new_n1708_), .ZN(new_n1712_));
  INV_X1    g1584(.A(new_n1706_), .ZN(new_n1713_));
  NAND2_X1  g1585(.A1(new_n1712_), .A2(new_n1713_), .ZN(new_n1714_));
  NAND3_X1  g1586(.A1(new_n1705_), .A2(new_n1706_), .A3(new_n1708_), .ZN(new_n1715_));
  OAI21_X1  g1587(.A(new_n1545_), .B1(new_n1540_), .B2(new_n1542_), .ZN(new_n1716_));
  NAND3_X1  g1588(.A1(new_n1714_), .A2(new_n1715_), .A3(new_n1716_), .ZN(new_n1717_));
  NAND2_X1  g1589(.A1(new_n1711_), .A2(new_n1717_), .ZN(new_n1718_));
  AOI21_X1  g1590(.A(new_n1549_), .B1(new_n1546_), .B2(new_n1547_), .ZN(new_n1719_));
  XNOR2_X1  g1591(.A(new_n1718_), .B(new_n1719_), .ZN(G6160gat));
  NOR3_X1   g1592(.A1(new_n1709_), .A2(new_n1710_), .A3(new_n1551_), .ZN(new_n1721_));
  NAND3_X1  g1593(.A1(new_n1548_), .A2(new_n1382_), .A3(new_n1388_), .ZN(new_n1722_));
  AOI21_X1  g1594(.A(new_n1721_), .B1(new_n1722_), .B2(new_n1711_), .ZN(new_n1723_));
  NOR2_X1   g1595(.A1(new_n165_), .A2(new_n1384_), .ZN(new_n1724_));
  NAND3_X1  g1596(.A1(new_n1666_), .A2(new_n1672_), .A3(new_n1674_), .ZN(new_n1725_));
  NAND2_X1  g1597(.A1(new_n1725_), .A2(new_n1672_), .ZN(new_n1726_));
  INV_X1    g1598(.A(new_n1726_), .ZN(new_n1727_));
  NAND2_X1  g1599(.A1(new_n1671_), .A2(new_n1661_), .ZN(new_n1728_));
  INV_X1    g1600(.A(new_n1728_), .ZN(new_n1729_));
  NOR2_X1   g1601(.A1(new_n377_), .A2(new_n648_), .ZN(new_n1730_));
  NOR2_X1   g1602(.A1(new_n542_), .A2(new_n533_), .ZN(new_n1731_));
  NOR2_X1   g1603(.A1(new_n1409_), .A2(new_n133_), .ZN(new_n1732_));
  OAI21_X1  g1604(.A(new_n1576_), .B1(new_n1579_), .B2(new_n1732_), .ZN(new_n1733_));
  OAI21_X1  g1605(.A(new_n1733_), .B1(new_n1232_), .B2(new_n159_), .ZN(new_n1734_));
  OAI21_X1  g1606(.A(new_n1734_), .B1(new_n159_), .B2(new_n1733_), .ZN(new_n1735_));
  NOR2_X1   g1607(.A1(new_n1578_), .A2(new_n198_), .ZN(new_n1736_));
  XOR2_X1   g1608(.A(new_n1735_), .B(new_n1736_), .Z(new_n1737_));
  OAI21_X1  g1609(.A(new_n1589_), .B1(new_n1586_), .B2(new_n1588_), .ZN(new_n1738_));
  AND2_X1   g1610(.A1(new_n1738_), .A2(new_n1572_), .ZN(new_n1739_));
  NOR2_X1   g1611(.A1(new_n1586_), .A2(new_n1582_), .ZN(new_n1740_));
  OAI21_X1  g1612(.A(new_n1737_), .B1(new_n1739_), .B2(new_n1740_), .ZN(new_n1741_));
  NAND2_X1  g1613(.A1(new_n1583_), .A2(new_n1572_), .ZN(new_n1742_));
  OAI21_X1  g1614(.A(new_n1742_), .B1(new_n1586_), .B2(new_n1582_), .ZN(new_n1743_));
  OR2_X1    g1615(.A1(new_n1743_), .A2(new_n1737_), .ZN(new_n1744_));
  NAND2_X1  g1616(.A1(new_n1741_), .A2(new_n1744_), .ZN(new_n1745_));
  NOR2_X1   g1617(.A1(new_n1406_), .A2(new_n276_), .ZN(new_n1746_));
  NAND2_X1  g1618(.A1(new_n1745_), .A2(new_n1746_), .ZN(new_n1747_));
  OAI211_X1 g1619(.A(new_n1741_), .B(new_n1744_), .C1(new_n1406_), .C2(new_n276_), .ZN(new_n1748_));
  NAND2_X1  g1620(.A1(new_n1603_), .A2(KEYINPUT48), .ZN(new_n1749_));
  NAND2_X1  g1621(.A1(new_n1749_), .A2(new_n1592_), .ZN(new_n1750_));
  NOR2_X1   g1622(.A1(new_n1603_), .A2(KEYINPUT48), .ZN(new_n1751_));
  OAI211_X1 g1623(.A(new_n1747_), .B(new_n1748_), .C1(new_n1750_), .C2(new_n1751_), .ZN(new_n1752_));
  NOR2_X1   g1624(.A1(new_n1260_), .A2(new_n289_), .ZN(new_n1753_));
  INV_X1    g1625(.A(new_n1753_), .ZN(new_n1754_));
  NAND2_X1  g1626(.A1(new_n1747_), .A2(new_n1748_), .ZN(new_n1755_));
  NAND3_X1  g1627(.A1(new_n1755_), .A2(new_n1592_), .A3(new_n1603_), .ZN(new_n1756_));
  NAND3_X1  g1628(.A1(new_n1752_), .A2(new_n1754_), .A3(new_n1756_), .ZN(new_n1757_));
  INV_X1    g1629(.A(new_n1757_), .ZN(new_n1758_));
  NAND2_X1  g1630(.A1(new_n1609_), .A2(new_n1607_), .ZN(new_n1759_));
  INV_X1    g1631(.A(new_n1759_), .ZN(new_n1760_));
  AOI21_X1  g1632(.A(new_n1754_), .B1(new_n1752_), .B2(new_n1756_), .ZN(new_n1761_));
  NOR3_X1   g1633(.A1(new_n1758_), .A2(new_n1760_), .A3(new_n1761_), .ZN(new_n1762_));
  INV_X1    g1634(.A(new_n1762_), .ZN(new_n1763_));
  OAI21_X1  g1635(.A(new_n1760_), .B1(new_n1758_), .B2(new_n1761_), .ZN(new_n1764_));
  OAI211_X1 g1636(.A(new_n1763_), .B(new_n1764_), .C1(new_n1084_), .C2(new_n363_), .ZN(new_n1765_));
  INV_X1    g1637(.A(new_n1764_), .ZN(new_n1766_));
  OAI211_X1 g1638(.A(G188gat), .B(G392gat), .C1(new_n1766_), .C2(new_n1762_), .ZN(new_n1767_));
  NAND2_X1  g1639(.A1(new_n1765_), .A2(new_n1767_), .ZN(new_n1768_));
  NAND2_X1  g1640(.A1(new_n1619_), .A2(KEYINPUT49), .ZN(new_n1769_));
  NAND3_X1  g1641(.A1(new_n1613_), .A2(new_n1616_), .A3(new_n1618_), .ZN(new_n1770_));
  INV_X1    g1642(.A(KEYINPUT49), .ZN(new_n1771_));
  AOI22_X1  g1643(.A1(new_n1770_), .A2(new_n1771_), .B1(new_n1612_), .B2(new_n1610_), .ZN(new_n1772_));
  AOI21_X1  g1644(.A(new_n1768_), .B1(new_n1769_), .B2(new_n1772_), .ZN(new_n1773_));
  INV_X1    g1645(.A(new_n1773_), .ZN(new_n1774_));
  NOR2_X1   g1646(.A1(new_n543_), .A2(new_n443_), .ZN(new_n1775_));
  NAND2_X1  g1647(.A1(new_n1775_), .A2(KEYINPUT50), .ZN(new_n1776_));
  NAND3_X1  g1648(.A1(new_n1768_), .A2(new_n1769_), .A3(new_n1772_), .ZN(new_n1777_));
  OR2_X1    g1649(.A1(new_n1775_), .A2(KEYINPUT50), .ZN(new_n1778_));
  NAND4_X1  g1650(.A1(new_n1774_), .A2(new_n1776_), .A3(new_n1777_), .A4(new_n1778_), .ZN(new_n1779_));
  NAND2_X1  g1651(.A1(new_n1630_), .A2(new_n1625_), .ZN(new_n1780_));
  INV_X1    g1652(.A(new_n1777_), .ZN(new_n1781_));
  OAI211_X1 g1653(.A(KEYINPUT50), .B(new_n1775_), .C1(new_n1781_), .C2(new_n1773_), .ZN(new_n1782_));
  NAND3_X1  g1654(.A1(new_n1779_), .A2(new_n1780_), .A3(new_n1782_), .ZN(new_n1783_));
  INV_X1    g1655(.A(new_n1783_), .ZN(new_n1784_));
  AOI21_X1  g1656(.A(new_n1780_), .B1(new_n1779_), .B2(new_n1782_), .ZN(new_n1785_));
  OAI21_X1  g1657(.A(new_n1731_), .B1(new_n1784_), .B2(new_n1785_), .ZN(new_n1786_));
  INV_X1    g1658(.A(new_n1785_), .ZN(new_n1787_));
  INV_X1    g1659(.A(new_n1731_), .ZN(new_n1788_));
  NAND3_X1  g1660(.A1(new_n1787_), .A2(new_n1788_), .A3(new_n1783_), .ZN(new_n1789_));
  NAND2_X1  g1661(.A1(new_n1643_), .A2(new_n1641_), .ZN(new_n1790_));
  NAND3_X1  g1662(.A1(new_n1786_), .A2(new_n1789_), .A3(new_n1790_), .ZN(new_n1791_));
  INV_X1    g1663(.A(new_n1791_), .ZN(new_n1792_));
  AOI21_X1  g1664(.A(new_n1790_), .B1(new_n1786_), .B2(new_n1789_), .ZN(new_n1793_));
  OAI21_X1  g1665(.A(new_n1730_), .B1(new_n1792_), .B2(new_n1793_), .ZN(new_n1794_));
  NAND2_X1  g1666(.A1(new_n1786_), .A2(new_n1789_), .ZN(new_n1795_));
  INV_X1    g1667(.A(new_n1790_), .ZN(new_n1796_));
  NAND2_X1  g1668(.A1(new_n1795_), .A2(new_n1796_), .ZN(new_n1797_));
  INV_X1    g1669(.A(new_n1730_), .ZN(new_n1798_));
  NAND3_X1  g1670(.A1(new_n1797_), .A2(new_n1798_), .A3(new_n1791_), .ZN(new_n1799_));
  AND2_X1   g1671(.A1(new_n1794_), .A2(new_n1799_), .ZN(new_n1800_));
  NAND2_X1  g1672(.A1(new_n1646_), .A2(new_n1650_), .ZN(new_n1801_));
  NAND2_X1  g1673(.A1(new_n1660_), .A2(new_n1801_), .ZN(new_n1802_));
  NAND2_X1  g1674(.A1(new_n1800_), .A2(new_n1802_), .ZN(new_n1803_));
  NOR2_X1   g1675(.A1(new_n300_), .A2(new_n654_), .ZN(new_n1804_));
  INV_X1    g1676(.A(new_n1804_), .ZN(new_n1805_));
  NAND2_X1  g1677(.A1(new_n1794_), .A2(new_n1799_), .ZN(new_n1806_));
  NAND3_X1  g1678(.A1(new_n1806_), .A2(new_n1660_), .A3(new_n1801_), .ZN(new_n1807_));
  NAND3_X1  g1679(.A1(new_n1803_), .A2(new_n1805_), .A3(new_n1807_), .ZN(new_n1808_));
  INV_X1    g1680(.A(new_n1808_), .ZN(new_n1809_));
  AOI21_X1  g1681(.A(new_n1805_), .B1(new_n1803_), .B2(new_n1807_), .ZN(new_n1810_));
  OAI21_X1  g1682(.A(new_n1729_), .B1(new_n1809_), .B2(new_n1810_), .ZN(new_n1811_));
  NAND2_X1  g1683(.A1(new_n1803_), .A2(new_n1807_), .ZN(new_n1812_));
  NAND2_X1  g1684(.A1(new_n1812_), .A2(new_n1804_), .ZN(new_n1813_));
  NAND3_X1  g1685(.A1(new_n1813_), .A2(new_n1728_), .A3(new_n1808_), .ZN(new_n1814_));
  NAND2_X1  g1686(.A1(G103gat), .A2(G477gat), .ZN(new_n1815_));
  AND3_X1   g1687(.A1(new_n1811_), .A2(new_n1814_), .A3(new_n1815_), .ZN(new_n1816_));
  AOI21_X1  g1688(.A(new_n1815_), .B1(new_n1811_), .B2(new_n1814_), .ZN(new_n1817_));
  OAI21_X1  g1689(.A(new_n1727_), .B1(new_n1816_), .B2(new_n1817_), .ZN(new_n1818_));
  NOR3_X1   g1690(.A1(new_n1809_), .A2(new_n1729_), .A3(new_n1810_), .ZN(new_n1819_));
  AOI21_X1  g1691(.A(new_n1728_), .B1(new_n1813_), .B2(new_n1808_), .ZN(new_n1820_));
  OAI211_X1 g1692(.A(G103gat), .B(G477gat), .C1(new_n1819_), .C2(new_n1820_), .ZN(new_n1821_));
  NAND3_X1  g1693(.A1(new_n1811_), .A2(new_n1814_), .A3(new_n1815_), .ZN(new_n1822_));
  NAND3_X1  g1694(.A1(new_n1821_), .A2(new_n1726_), .A3(new_n1822_), .ZN(new_n1823_));
  NAND2_X1  g1695(.A1(G86gat), .A2(G494gat), .ZN(new_n1824_));
  AND3_X1   g1696(.A1(new_n1818_), .A2(new_n1823_), .A3(new_n1824_), .ZN(new_n1825_));
  AOI21_X1  g1697(.A(new_n1824_), .B1(new_n1818_), .B2(new_n1823_), .ZN(new_n1826_));
  OAI211_X1 g1698(.A(new_n1684_), .B(new_n1680_), .C1(new_n1825_), .C2(new_n1826_), .ZN(new_n1827_));
  NAND2_X1  g1699(.A1(new_n1818_), .A2(new_n1823_), .ZN(new_n1828_));
  NAND3_X1  g1700(.A1(new_n1828_), .A2(G86gat), .A3(G494gat), .ZN(new_n1829_));
  NAND2_X1  g1701(.A1(new_n1684_), .A2(new_n1680_), .ZN(new_n1830_));
  NAND3_X1  g1702(.A1(new_n1818_), .A2(new_n1823_), .A3(new_n1824_), .ZN(new_n1831_));
  NAND3_X1  g1703(.A1(new_n1829_), .A2(new_n1830_), .A3(new_n1831_), .ZN(new_n1832_));
  NAND2_X1  g1704(.A1(new_n1827_), .A2(new_n1832_), .ZN(new_n1833_));
  NOR2_X1   g1705(.A1(new_n166_), .A2(new_n1218_), .ZN(new_n1834_));
  NAND2_X1  g1706(.A1(new_n1833_), .A2(new_n1834_), .ZN(new_n1835_));
  INV_X1    g1707(.A(new_n1834_), .ZN(new_n1836_));
  NAND3_X1  g1708(.A1(new_n1827_), .A2(new_n1832_), .A3(new_n1836_), .ZN(new_n1837_));
  NAND2_X1  g1709(.A1(new_n1688_), .A2(new_n1689_), .ZN(new_n1838_));
  AOI22_X1  g1710(.A1(new_n1835_), .A2(new_n1837_), .B1(new_n1693_), .B2(new_n1838_), .ZN(new_n1839_));
  AND3_X1   g1711(.A1(new_n1827_), .A2(new_n1832_), .A3(new_n1836_), .ZN(new_n1840_));
  AOI21_X1  g1712(.A(new_n1836_), .B1(new_n1827_), .B2(new_n1832_), .ZN(new_n1841_));
  NAND2_X1  g1713(.A1(new_n1838_), .A2(new_n1693_), .ZN(new_n1842_));
  NOR3_X1   g1714(.A1(new_n1840_), .A2(new_n1841_), .A3(new_n1842_), .ZN(new_n1843_));
  OAI21_X1  g1715(.A(new_n1724_), .B1(new_n1839_), .B2(new_n1843_), .ZN(new_n1844_));
  OAI21_X1  g1716(.A(new_n1842_), .B1(new_n1840_), .B2(new_n1841_), .ZN(new_n1845_));
  NAND4_X1  g1717(.A1(new_n1835_), .A2(new_n1693_), .A3(new_n1837_), .A4(new_n1838_), .ZN(new_n1846_));
  OAI211_X1 g1718(.A(new_n1845_), .B(new_n1846_), .C1(new_n165_), .C2(new_n1384_), .ZN(new_n1847_));
  NAND2_X1  g1719(.A1(new_n1844_), .A2(new_n1847_), .ZN(new_n1848_));
  NAND2_X1  g1720(.A1(new_n1701_), .A2(new_n1703_), .ZN(new_n1849_));
  NAND3_X1  g1721(.A1(new_n1848_), .A2(new_n1714_), .A3(new_n1849_), .ZN(new_n1850_));
  INV_X1    g1722(.A(new_n1849_), .ZN(new_n1851_));
  OAI211_X1 g1723(.A(new_n1847_), .B(new_n1844_), .C1(new_n1710_), .C2(new_n1851_), .ZN(new_n1852_));
  NAND2_X1  g1724(.A1(new_n1850_), .A2(new_n1852_), .ZN(new_n1853_));
  XNOR2_X1  g1725(.A(new_n1723_), .B(new_n1853_), .ZN(G6170gat));
  OAI21_X1  g1726(.A(new_n1852_), .B1(new_n1723_), .B2(new_n1853_), .ZN(new_n1855_));
  NAND2_X1  g1727(.A1(G86gat), .A2(G511gat), .ZN(new_n1856_));
  NAND2_X1  g1728(.A1(G103gat), .A2(G494gat), .ZN(new_n1857_));
  NAND2_X1  g1729(.A1(G137gat), .A2(G460gat), .ZN(new_n1858_));
  NAND2_X1  g1730(.A1(G171gat), .A2(G426gat), .ZN(new_n1859_));
  XOR2_X1   g1731(.A(new_n1859_), .B(KEYINPUT51), .Z(new_n1860_));
  INV_X1    g1732(.A(new_n1860_), .ZN(new_n1861_));
  AND2_X1   g1733(.A1(new_n1757_), .A2(new_n1752_), .ZN(new_n1862_));
  OAI21_X1  g1734(.A(new_n1734_), .B1(new_n1735_), .B2(new_n1736_), .ZN(new_n1863_));
  NAND2_X1  g1735(.A1(G256gat), .A2(G341gat), .ZN(new_n1864_));
  XNOR2_X1  g1736(.A(new_n1863_), .B(new_n1864_), .ZN(new_n1865_));
  NOR2_X1   g1737(.A1(new_n1578_), .A2(new_n276_), .ZN(new_n1866_));
  XNOR2_X1  g1738(.A(new_n1865_), .B(new_n1866_), .ZN(new_n1867_));
  NAND2_X1  g1739(.A1(new_n1743_), .A2(new_n1737_), .ZN(new_n1868_));
  NAND2_X1  g1740(.A1(new_n1868_), .A2(new_n1746_), .ZN(new_n1869_));
  NAND2_X1  g1741(.A1(new_n1869_), .A2(new_n1744_), .ZN(new_n1870_));
  XNOR2_X1  g1742(.A(new_n1867_), .B(new_n1870_), .ZN(new_n1871_));
  NOR2_X1   g1743(.A1(new_n1406_), .A2(new_n289_), .ZN(new_n1872_));
  XNOR2_X1  g1744(.A(new_n1871_), .B(new_n1872_), .ZN(new_n1873_));
  OR2_X1    g1745(.A1(new_n1862_), .A2(new_n1873_), .ZN(new_n1874_));
  NAND2_X1  g1746(.A1(new_n1862_), .A2(new_n1873_), .ZN(new_n1875_));
  NAND2_X1  g1747(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1876_));
  NAND3_X1  g1748(.A1(new_n1876_), .A2(G205gat), .A3(G392gat), .ZN(new_n1877_));
  OAI211_X1 g1749(.A(new_n1874_), .B(new_n1875_), .C1(new_n1260_), .C2(new_n363_), .ZN(new_n1878_));
  NAND2_X1  g1750(.A1(new_n1877_), .A2(new_n1878_), .ZN(new_n1879_));
  NAND3_X1  g1751(.A1(new_n1879_), .A2(new_n1763_), .A3(new_n1765_), .ZN(new_n1880_));
  NOR2_X1   g1752(.A1(new_n1084_), .A2(new_n443_), .ZN(new_n1881_));
  INV_X1    g1753(.A(new_n1881_), .ZN(new_n1882_));
  NAND2_X1  g1754(.A1(new_n1765_), .A2(new_n1763_), .ZN(new_n1883_));
  NAND3_X1  g1755(.A1(new_n1883_), .A2(new_n1878_), .A3(new_n1877_), .ZN(new_n1884_));
  NAND3_X1  g1756(.A1(new_n1880_), .A2(new_n1882_), .A3(new_n1884_), .ZN(new_n1885_));
  INV_X1    g1757(.A(new_n1885_), .ZN(new_n1886_));
  AOI21_X1  g1758(.A(new_n1882_), .B1(new_n1880_), .B2(new_n1884_), .ZN(new_n1887_));
  NOR2_X1   g1759(.A1(new_n1886_), .A2(new_n1887_), .ZN(new_n1888_));
  OAI21_X1  g1760(.A(new_n1777_), .B1(new_n543_), .B2(new_n443_), .ZN(new_n1889_));
  NAND2_X1  g1761(.A1(new_n1889_), .A2(new_n1774_), .ZN(new_n1890_));
  NAND2_X1  g1762(.A1(new_n1888_), .A2(new_n1890_), .ZN(new_n1891_));
  INV_X1    g1763(.A(new_n1891_), .ZN(new_n1892_));
  NOR2_X1   g1764(.A1(new_n1888_), .A2(new_n1890_), .ZN(new_n1893_));
  OAI21_X1  g1765(.A(new_n1861_), .B1(new_n1892_), .B2(new_n1893_), .ZN(new_n1894_));
  OR2_X1    g1766(.A1(new_n1888_), .A2(new_n1890_), .ZN(new_n1895_));
  NAND3_X1  g1767(.A1(new_n1895_), .A2(new_n1860_), .A3(new_n1891_), .ZN(new_n1896_));
  NAND2_X1  g1768(.A1(new_n1894_), .A2(new_n1896_), .ZN(new_n1897_));
  NAND2_X1  g1769(.A1(new_n1789_), .A2(new_n1783_), .ZN(new_n1898_));
  INV_X1    g1770(.A(new_n1898_), .ZN(new_n1899_));
  NAND2_X1  g1771(.A1(new_n1897_), .A2(new_n1899_), .ZN(new_n1900_));
  NAND2_X1  g1772(.A1(G154gat), .A2(G443gat), .ZN(new_n1901_));
  NAND3_X1  g1773(.A1(new_n1898_), .A2(new_n1894_), .A3(new_n1896_), .ZN(new_n1902_));
  AND3_X1   g1774(.A1(new_n1900_), .A2(new_n1901_), .A3(new_n1902_), .ZN(new_n1903_));
  AOI21_X1  g1775(.A(new_n1901_), .B1(new_n1900_), .B2(new_n1902_), .ZN(new_n1904_));
  OAI211_X1 g1776(.A(new_n1791_), .B(new_n1799_), .C1(new_n1903_), .C2(new_n1904_), .ZN(new_n1905_));
  INV_X1    g1777(.A(new_n1904_), .ZN(new_n1906_));
  NAND2_X1  g1778(.A1(new_n1799_), .A2(new_n1791_), .ZN(new_n1907_));
  NAND3_X1  g1779(.A1(new_n1900_), .A2(new_n1901_), .A3(new_n1902_), .ZN(new_n1908_));
  NAND3_X1  g1780(.A1(new_n1906_), .A2(new_n1907_), .A3(new_n1908_), .ZN(new_n1909_));
  AOI21_X1  g1781(.A(new_n1858_), .B1(new_n1905_), .B2(new_n1909_), .ZN(new_n1910_));
  INV_X1    g1782(.A(new_n1910_), .ZN(new_n1911_));
  NAND3_X1  g1783(.A1(new_n1905_), .A2(new_n1909_), .A3(new_n1858_), .ZN(new_n1912_));
  NAND2_X1  g1784(.A1(new_n1911_), .A2(new_n1912_), .ZN(new_n1913_));
  NAND2_X1  g1785(.A1(new_n1808_), .A2(new_n1803_), .ZN(new_n1914_));
  INV_X1    g1786(.A(new_n1914_), .ZN(new_n1915_));
  NAND2_X1  g1787(.A1(new_n1913_), .A2(new_n1915_), .ZN(new_n1916_));
  NAND3_X1  g1788(.A1(new_n1911_), .A2(new_n1914_), .A3(new_n1912_), .ZN(new_n1917_));
  NAND2_X1  g1789(.A1(new_n1916_), .A2(new_n1917_), .ZN(new_n1918_));
  NOR2_X1   g1790(.A1(new_n300_), .A2(new_n890_), .ZN(new_n1919_));
  NAND2_X1  g1791(.A1(new_n1918_), .A2(new_n1919_), .ZN(new_n1920_));
  OAI211_X1 g1792(.A(new_n1916_), .B(new_n1917_), .C1(new_n300_), .C2(new_n890_), .ZN(new_n1921_));
  NAND2_X1  g1793(.A1(new_n1920_), .A2(new_n1921_), .ZN(new_n1922_));
  NOR2_X1   g1794(.A1(new_n1816_), .A2(new_n1819_), .ZN(new_n1923_));
  NAND2_X1  g1795(.A1(new_n1922_), .A2(new_n1923_), .ZN(new_n1924_));
  OAI211_X1 g1796(.A(new_n1920_), .B(new_n1921_), .C1(new_n1819_), .C2(new_n1816_), .ZN(new_n1925_));
  AOI21_X1  g1797(.A(new_n1857_), .B1(new_n1924_), .B2(new_n1925_), .ZN(new_n1926_));
  INV_X1    g1798(.A(new_n1926_), .ZN(new_n1927_));
  NAND2_X1  g1799(.A1(new_n1831_), .A2(new_n1823_), .ZN(new_n1928_));
  NAND3_X1  g1800(.A1(new_n1924_), .A2(new_n1857_), .A3(new_n1925_), .ZN(new_n1929_));
  NAND3_X1  g1801(.A1(new_n1927_), .A2(new_n1928_), .A3(new_n1929_), .ZN(new_n1930_));
  INV_X1    g1802(.A(new_n1928_), .ZN(new_n1931_));
  AND3_X1   g1803(.A1(new_n1924_), .A2(new_n1857_), .A3(new_n1925_), .ZN(new_n1932_));
  OAI21_X1  g1804(.A(new_n1931_), .B1(new_n1932_), .B2(new_n1926_), .ZN(new_n1933_));
  AOI21_X1  g1805(.A(new_n1856_), .B1(new_n1930_), .B2(new_n1933_), .ZN(new_n1934_));
  INV_X1    g1806(.A(new_n1934_), .ZN(new_n1935_));
  NAND2_X1  g1807(.A1(new_n1837_), .A2(new_n1832_), .ZN(new_n1936_));
  NAND3_X1  g1808(.A1(new_n1930_), .A2(new_n1933_), .A3(new_n1856_), .ZN(new_n1937_));
  NAND3_X1  g1809(.A1(new_n1935_), .A2(new_n1936_), .A3(new_n1937_), .ZN(new_n1938_));
  INV_X1    g1810(.A(new_n1936_), .ZN(new_n1939_));
  AND3_X1   g1811(.A1(new_n1930_), .A2(new_n1856_), .A3(new_n1933_), .ZN(new_n1940_));
  OAI21_X1  g1812(.A(new_n1939_), .B1(new_n1940_), .B2(new_n1934_), .ZN(new_n1941_));
  NAND2_X1  g1813(.A1(new_n1938_), .A2(new_n1941_), .ZN(new_n1942_));
  NAND3_X1  g1814(.A1(new_n1942_), .A2(G69gat), .A3(G528gat), .ZN(new_n1943_));
  NAND2_X1  g1815(.A1(new_n1847_), .A2(new_n1846_), .ZN(new_n1944_));
  OAI211_X1 g1816(.A(new_n1938_), .B(new_n1941_), .C1(new_n166_), .C2(new_n1384_), .ZN(new_n1945_));
  AND3_X1   g1817(.A1(new_n1943_), .A2(new_n1944_), .A3(new_n1945_), .ZN(new_n1946_));
  AOI21_X1  g1818(.A(new_n1944_), .B1(new_n1943_), .B2(new_n1945_), .ZN(new_n1947_));
  NOR2_X1   g1819(.A1(new_n1946_), .A2(new_n1947_), .ZN(new_n1948_));
  XNOR2_X1  g1820(.A(new_n1855_), .B(new_n1948_), .ZN(G6180gat));
  INV_X1    g1821(.A(new_n1946_), .ZN(new_n1950_));
  INV_X1    g1822(.A(new_n1852_), .ZN(new_n1951_));
  AOI21_X1  g1823(.A(new_n1716_), .B1(new_n1714_), .B2(new_n1715_), .ZN(new_n1952_));
  OAI21_X1  g1824(.A(new_n1717_), .B1(new_n1952_), .B2(new_n1719_), .ZN(new_n1953_));
  AOI21_X1  g1825(.A(new_n1951_), .B1(new_n1953_), .B2(new_n1850_), .ZN(new_n1954_));
  OAI21_X1  g1826(.A(new_n1950_), .B1(new_n1954_), .B2(new_n1947_), .ZN(new_n1955_));
  NAND2_X1  g1827(.A1(new_n1937_), .A2(new_n1930_), .ZN(new_n1956_));
  INV_X1    g1828(.A(new_n1956_), .ZN(new_n1957_));
  NAND2_X1  g1829(.A1(new_n1929_), .A2(new_n1925_), .ZN(new_n1958_));
  INV_X1    g1830(.A(new_n1958_), .ZN(new_n1959_));
  XNOR2_X1  g1831(.A(new_n1902_), .B(KEYINPUT53), .ZN(new_n1960_));
  NAND2_X1  g1832(.A1(new_n1960_), .A2(new_n1908_), .ZN(new_n1961_));
  INV_X1    g1833(.A(new_n1961_), .ZN(new_n1962_));
  INV_X1    g1834(.A(KEYINPUT54), .ZN(new_n1963_));
  NOR2_X1   g1835(.A1(new_n1865_), .A2(new_n1866_), .ZN(new_n1964_));
  AOI21_X1  g1836(.A(new_n1964_), .B1(new_n1863_), .B2(new_n1864_), .ZN(new_n1965_));
  NOR2_X1   g1837(.A1(new_n1232_), .A2(new_n276_), .ZN(new_n1966_));
  INV_X1    g1838(.A(new_n1966_), .ZN(new_n1967_));
  NOR2_X1   g1839(.A1(new_n1967_), .A2(KEYINPUT52), .ZN(new_n1968_));
  INV_X1    g1840(.A(KEYINPUT52), .ZN(new_n1969_));
  NOR2_X1   g1841(.A1(new_n1966_), .A2(new_n1969_), .ZN(new_n1970_));
  OAI21_X1  g1842(.A(new_n1965_), .B1(new_n1968_), .B2(new_n1970_), .ZN(new_n1971_));
  OAI21_X1  g1843(.A(new_n1971_), .B1(new_n1965_), .B2(new_n1970_), .ZN(new_n1972_));
  INV_X1    g1844(.A(new_n1972_), .ZN(new_n1973_));
  NOR2_X1   g1845(.A1(new_n1578_), .A2(new_n289_), .ZN(new_n1974_));
  NAND2_X1  g1846(.A1(new_n1973_), .A2(new_n1974_), .ZN(new_n1975_));
  INV_X1    g1847(.A(new_n1974_), .ZN(new_n1976_));
  NAND2_X1  g1848(.A1(new_n1972_), .A2(new_n1976_), .ZN(new_n1977_));
  NAND2_X1  g1849(.A1(new_n1975_), .A2(new_n1977_), .ZN(new_n1978_));
  OR2_X1    g1850(.A1(new_n1871_), .A2(new_n1872_), .ZN(new_n1979_));
  OR2_X1    g1851(.A1(new_n1867_), .A2(new_n1870_), .ZN(new_n1980_));
  NAND2_X1  g1852(.A1(new_n1979_), .A2(new_n1980_), .ZN(new_n1981_));
  XOR2_X1   g1853(.A(new_n1978_), .B(new_n1981_), .Z(new_n1982_));
  NOR2_X1   g1854(.A1(new_n1406_), .A2(new_n363_), .ZN(new_n1983_));
  XNOR2_X1  g1855(.A(new_n1982_), .B(new_n1983_), .ZN(new_n1984_));
  INV_X1    g1856(.A(new_n1984_), .ZN(new_n1985_));
  NAND2_X1  g1857(.A1(new_n1878_), .A2(new_n1874_), .ZN(new_n1986_));
  NAND2_X1  g1858(.A1(new_n1985_), .A2(new_n1986_), .ZN(new_n1987_));
  NAND3_X1  g1859(.A1(new_n1984_), .A2(new_n1874_), .A3(new_n1878_), .ZN(new_n1988_));
  NAND2_X1  g1860(.A1(new_n1987_), .A2(new_n1988_), .ZN(new_n1989_));
  NOR2_X1   g1861(.A1(new_n1260_), .A2(new_n443_), .ZN(new_n1990_));
  NAND2_X1  g1862(.A1(new_n1989_), .A2(new_n1990_), .ZN(new_n1991_));
  OAI211_X1 g1863(.A(new_n1987_), .B(new_n1988_), .C1(new_n1260_), .C2(new_n443_), .ZN(new_n1992_));
  NAND2_X1  g1864(.A1(new_n1991_), .A2(new_n1992_), .ZN(new_n1993_));
  NAND3_X1  g1865(.A1(new_n1993_), .A2(new_n1884_), .A3(new_n1885_), .ZN(new_n1994_));
  NAND2_X1  g1866(.A1(new_n1885_), .A2(new_n1884_), .ZN(new_n1995_));
  NAND3_X1  g1867(.A1(new_n1995_), .A2(new_n1992_), .A3(new_n1991_), .ZN(new_n1996_));
  NAND2_X1  g1868(.A1(new_n1994_), .A2(new_n1996_), .ZN(new_n1997_));
  NAND2_X1  g1869(.A1(G188gat), .A2(G426gat), .ZN(new_n1998_));
  XNOR2_X1  g1870(.A(new_n1997_), .B(new_n1998_), .ZN(new_n1999_));
  NAND2_X1  g1871(.A1(new_n1896_), .A2(new_n1891_), .ZN(new_n2000_));
  OR2_X1    g1872(.A1(new_n1999_), .A2(new_n2000_), .ZN(new_n2001_));
  NOR2_X1   g1873(.A1(new_n543_), .A2(new_n648_), .ZN(new_n2002_));
  INV_X1    g1874(.A(new_n2002_), .ZN(new_n2003_));
  NAND2_X1  g1875(.A1(new_n1999_), .A2(new_n2000_), .ZN(new_n2004_));
  NAND3_X1  g1876(.A1(new_n2001_), .A2(new_n2003_), .A3(new_n2004_), .ZN(new_n2005_));
  INV_X1    g1877(.A(new_n2005_), .ZN(new_n2006_));
  AOI21_X1  g1878(.A(new_n2003_), .B1(new_n2001_), .B2(new_n2004_), .ZN(new_n2007_));
  OAI21_X1  g1879(.A(new_n1963_), .B1(new_n2006_), .B2(new_n2007_), .ZN(new_n2008_));
  XNOR2_X1  g1880(.A(new_n1999_), .B(new_n2000_), .ZN(new_n2009_));
  NAND2_X1  g1881(.A1(new_n2009_), .A2(new_n2002_), .ZN(new_n2010_));
  NAND3_X1  g1882(.A1(new_n2010_), .A2(new_n2005_), .A3(KEYINPUT54), .ZN(new_n2011_));
  AOI21_X1  g1883(.A(new_n1962_), .B1(new_n2008_), .B2(new_n2011_), .ZN(new_n2012_));
  AOI21_X1  g1884(.A(KEYINPUT54), .B1(new_n2010_), .B2(new_n2005_), .ZN(new_n2013_));
  NOR2_X1   g1885(.A1(new_n2013_), .A2(new_n1961_), .ZN(new_n2014_));
  OAI22_X1  g1886(.A1(new_n2012_), .A2(new_n2014_), .B1(new_n542_), .B2(new_n654_), .ZN(new_n2015_));
  NOR3_X1   g1887(.A1(new_n2006_), .A2(new_n1963_), .A3(new_n2007_), .ZN(new_n2016_));
  OAI21_X1  g1888(.A(new_n1961_), .B1(new_n2016_), .B2(new_n2013_), .ZN(new_n2017_));
  NOR2_X1   g1889(.A1(new_n542_), .A2(new_n654_), .ZN(new_n2018_));
  NAND2_X1  g1890(.A1(new_n2008_), .A2(new_n1962_), .ZN(new_n2019_));
  NAND3_X1  g1891(.A1(new_n2017_), .A2(new_n2018_), .A3(new_n2019_), .ZN(new_n2020_));
  NAND2_X1  g1892(.A1(new_n2015_), .A2(new_n2020_), .ZN(new_n2021_));
  NAND2_X1  g1893(.A1(new_n1912_), .A2(new_n1909_), .ZN(new_n2022_));
  INV_X1    g1894(.A(new_n2022_), .ZN(new_n2023_));
  NAND2_X1  g1895(.A1(new_n2021_), .A2(new_n2023_), .ZN(new_n2024_));
  NAND2_X1  g1896(.A1(G137gat), .A2(G477gat), .ZN(new_n2025_));
  NAND3_X1  g1897(.A1(new_n2015_), .A2(new_n2020_), .A3(new_n2022_), .ZN(new_n2026_));
  AND3_X1   g1898(.A1(new_n2024_), .A2(new_n2025_), .A3(new_n2026_), .ZN(new_n2027_));
  AOI21_X1  g1899(.A(new_n2025_), .B1(new_n2024_), .B2(new_n2026_), .ZN(new_n2028_));
  OAI211_X1 g1900(.A(new_n1917_), .B(new_n1921_), .C1(new_n2027_), .C2(new_n2028_), .ZN(new_n2029_));
  INV_X1    g1901(.A(new_n2026_), .ZN(new_n2030_));
  AOI21_X1  g1902(.A(new_n2022_), .B1(new_n2015_), .B2(new_n2020_), .ZN(new_n2031_));
  OAI211_X1 g1903(.A(G137gat), .B(G477gat), .C1(new_n2030_), .C2(new_n2031_), .ZN(new_n2032_));
  NAND3_X1  g1904(.A1(new_n2024_), .A2(new_n2025_), .A3(new_n2026_), .ZN(new_n2033_));
  NAND2_X1  g1905(.A1(new_n1921_), .A2(new_n1917_), .ZN(new_n2034_));
  NAND3_X1  g1906(.A1(new_n2032_), .A2(new_n2033_), .A3(new_n2034_), .ZN(new_n2035_));
  NOR2_X1   g1907(.A1(new_n300_), .A2(new_n1057_), .ZN(new_n2036_));
  INV_X1    g1908(.A(new_n2036_), .ZN(new_n2037_));
  AND3_X1   g1909(.A1(new_n2029_), .A2(new_n2035_), .A3(new_n2037_), .ZN(new_n2038_));
  AOI21_X1  g1910(.A(new_n2037_), .B1(new_n2029_), .B2(new_n2035_), .ZN(new_n2039_));
  OAI21_X1  g1911(.A(new_n1959_), .B1(new_n2038_), .B2(new_n2039_), .ZN(new_n2040_));
  NAND2_X1  g1912(.A1(new_n2029_), .A2(new_n2035_), .ZN(new_n2041_));
  NAND2_X1  g1913(.A1(new_n2041_), .A2(new_n2036_), .ZN(new_n2042_));
  NAND3_X1  g1914(.A1(new_n2029_), .A2(new_n2035_), .A3(new_n2037_), .ZN(new_n2043_));
  NAND3_X1  g1915(.A1(new_n2042_), .A2(new_n1958_), .A3(new_n2043_), .ZN(new_n2044_));
  NOR2_X1   g1916(.A1(new_n243_), .A2(new_n1218_), .ZN(new_n2045_));
  INV_X1    g1917(.A(new_n2045_), .ZN(new_n2046_));
  NAND3_X1  g1918(.A1(new_n2040_), .A2(new_n2044_), .A3(new_n2046_), .ZN(new_n2047_));
  INV_X1    g1919(.A(new_n2047_), .ZN(new_n2048_));
  AOI21_X1  g1920(.A(new_n2046_), .B1(new_n2040_), .B2(new_n2044_), .ZN(new_n2049_));
  OAI21_X1  g1921(.A(new_n1957_), .B1(new_n2048_), .B2(new_n2049_), .ZN(new_n2050_));
  NAND2_X1  g1922(.A1(new_n2040_), .A2(new_n2044_), .ZN(new_n2051_));
  NAND2_X1  g1923(.A1(new_n2051_), .A2(new_n2045_), .ZN(new_n2052_));
  NAND3_X1  g1924(.A1(new_n2052_), .A2(new_n1956_), .A3(new_n2047_), .ZN(new_n2053_));
  NAND2_X1  g1925(.A1(new_n2050_), .A2(new_n2053_), .ZN(new_n2054_));
  NOR2_X1   g1926(.A1(new_n242_), .A2(new_n1384_), .ZN(new_n2055_));
  NAND2_X1  g1927(.A1(new_n2054_), .A2(new_n2055_), .ZN(new_n2056_));
  OAI211_X1 g1928(.A(new_n2050_), .B(new_n2053_), .C1(new_n242_), .C2(new_n1384_), .ZN(new_n2057_));
  NAND2_X1  g1929(.A1(new_n2056_), .A2(new_n2057_), .ZN(new_n2058_));
  NAND2_X1  g1930(.A1(new_n1945_), .A2(new_n1938_), .ZN(new_n2059_));
  XNOR2_X1  g1931(.A(new_n2058_), .B(new_n2059_), .ZN(new_n2060_));
  XNOR2_X1  g1932(.A(new_n1955_), .B(new_n2060_), .ZN(G6190gat));
  AOI21_X1  g1933(.A(new_n2058_), .B1(new_n1938_), .B2(new_n1945_), .ZN(new_n2062_));
  INV_X1    g1934(.A(new_n2062_), .ZN(new_n2063_));
  AOI21_X1  g1935(.A(new_n1946_), .B1(new_n1855_), .B2(new_n1948_), .ZN(new_n2064_));
  AOI21_X1  g1936(.A(new_n2059_), .B1(new_n2056_), .B2(new_n2057_), .ZN(new_n2065_));
  OAI21_X1  g1937(.A(new_n2063_), .B1(new_n2064_), .B2(new_n2065_), .ZN(new_n2066_));
  NAND2_X1  g1938(.A1(G137gat), .A2(G494gat), .ZN(new_n2067_));
  NOR2_X1   g1939(.A1(new_n542_), .A2(new_n890_), .ZN(new_n2068_));
  OAI21_X1  g1940(.A(new_n1977_), .B1(new_n1965_), .B2(new_n1966_), .ZN(new_n2069_));
  NOR2_X1   g1941(.A1(new_n1232_), .A2(new_n289_), .ZN(new_n2070_));
  XNOR2_X1  g1942(.A(new_n2069_), .B(new_n2070_), .ZN(new_n2071_));
  NAND2_X1  g1943(.A1(G239gat), .A2(G392gat), .ZN(new_n2072_));
  XOR2_X1   g1944(.A(new_n2072_), .B(KEYINPUT55), .Z(new_n2073_));
  NAND2_X1  g1945(.A1(new_n2071_), .A2(new_n2073_), .ZN(new_n2074_));
  OR2_X1    g1946(.A1(new_n2074_), .A2(KEYINPUT56), .ZN(new_n2075_));
  INV_X1    g1947(.A(new_n2071_), .ZN(new_n2076_));
  NAND2_X1  g1948(.A1(new_n2076_), .A2(new_n2072_), .ZN(new_n2077_));
  NAND2_X1  g1949(.A1(new_n2074_), .A2(KEYINPUT56), .ZN(new_n2078_));
  NAND3_X1  g1950(.A1(new_n2075_), .A2(new_n2077_), .A3(new_n2078_), .ZN(new_n2079_));
  NAND3_X1  g1951(.A1(new_n1981_), .A2(new_n1975_), .A3(new_n1977_), .ZN(new_n2080_));
  OAI21_X1  g1952(.A(new_n2080_), .B1(new_n1982_), .B2(new_n1983_), .ZN(new_n2081_));
  XNOR2_X1  g1953(.A(new_n2079_), .B(new_n2081_), .ZN(new_n2082_));
  NOR2_X1   g1954(.A1(new_n1406_), .A2(new_n443_), .ZN(new_n2083_));
  XNOR2_X1  g1955(.A(new_n2082_), .B(new_n2083_), .ZN(new_n2084_));
  AND2_X1   g1956(.A1(new_n1992_), .A2(new_n1987_), .ZN(new_n2085_));
  OR2_X1    g1957(.A1(new_n2084_), .A2(new_n2085_), .ZN(new_n2086_));
  NAND2_X1  g1958(.A1(new_n2084_), .A2(new_n2085_), .ZN(new_n2087_));
  NAND2_X1  g1959(.A1(new_n2086_), .A2(new_n2087_), .ZN(new_n2088_));
  NOR2_X1   g1960(.A1(new_n1260_), .A2(new_n533_), .ZN(new_n2089_));
  NAND2_X1  g1961(.A1(new_n2088_), .A2(new_n2089_), .ZN(new_n2090_));
  XOR2_X1   g1962(.A(new_n2089_), .B(KEYINPUT57), .Z(new_n2091_));
  NAND3_X1  g1963(.A1(new_n2086_), .A2(new_n2087_), .A3(new_n2091_), .ZN(new_n2092_));
  NAND2_X1  g1964(.A1(new_n2090_), .A2(new_n2092_), .ZN(new_n2093_));
  NAND3_X1  g1965(.A1(new_n1994_), .A2(new_n1998_), .A3(new_n1996_), .ZN(new_n2094_));
  NAND3_X1  g1966(.A1(new_n2093_), .A2(new_n1996_), .A3(new_n2094_), .ZN(new_n2095_));
  NAND2_X1  g1967(.A1(G188gat), .A2(G443gat), .ZN(new_n2096_));
  NAND2_X1  g1968(.A1(new_n2094_), .A2(new_n1996_), .ZN(new_n2097_));
  NAND3_X1  g1969(.A1(new_n2090_), .A2(new_n2097_), .A3(new_n2092_), .ZN(new_n2098_));
  NAND3_X1  g1970(.A1(new_n2095_), .A2(new_n2096_), .A3(new_n2098_), .ZN(new_n2099_));
  INV_X1    g1971(.A(new_n2099_), .ZN(new_n2100_));
  AOI21_X1  g1972(.A(new_n2096_), .B1(new_n2095_), .B2(new_n2098_), .ZN(new_n2101_));
  NOR2_X1   g1973(.A1(new_n2100_), .A2(new_n2101_), .ZN(new_n2102_));
  NAND2_X1  g1974(.A1(new_n2005_), .A2(new_n2004_), .ZN(new_n2103_));
  OR2_X1    g1975(.A1(new_n2102_), .A2(new_n2103_), .ZN(new_n2104_));
  NAND2_X1  g1976(.A1(new_n2102_), .A2(new_n2103_), .ZN(new_n2105_));
  NAND2_X1  g1977(.A1(new_n2104_), .A2(new_n2105_), .ZN(new_n2106_));
  NAND3_X1  g1978(.A1(new_n2106_), .A2(G171gat), .A3(G460gat), .ZN(new_n2107_));
  OAI211_X1 g1979(.A(new_n2104_), .B(new_n2105_), .C1(new_n543_), .C2(new_n654_), .ZN(new_n2108_));
  NAND2_X1  g1980(.A1(new_n2107_), .A2(new_n2108_), .ZN(new_n2109_));
  NAND3_X1  g1981(.A1(new_n2010_), .A2(new_n1961_), .A3(new_n2005_), .ZN(new_n2110_));
  AND2_X1   g1982(.A1(new_n2015_), .A2(new_n2110_), .ZN(new_n2111_));
  NAND2_X1  g1983(.A1(new_n2109_), .A2(new_n2111_), .ZN(new_n2112_));
  INV_X1    g1984(.A(new_n2112_), .ZN(new_n2113_));
  NOR2_X1   g1985(.A1(new_n2109_), .A2(new_n2111_), .ZN(new_n2114_));
  OAI21_X1  g1986(.A(new_n2068_), .B1(new_n2113_), .B2(new_n2114_), .ZN(new_n2115_));
  INV_X1    g1987(.A(new_n2114_), .ZN(new_n2116_));
  INV_X1    g1988(.A(new_n2068_), .ZN(new_n2117_));
  NAND3_X1  g1989(.A1(new_n2116_), .A2(new_n2117_), .A3(new_n2112_), .ZN(new_n2118_));
  NAND2_X1  g1990(.A1(new_n2115_), .A2(new_n2118_), .ZN(new_n2119_));
  NAND2_X1  g1991(.A1(new_n2033_), .A2(new_n2026_), .ZN(new_n2120_));
  INV_X1    g1992(.A(new_n2120_), .ZN(new_n2121_));
  NAND2_X1  g1993(.A1(new_n2119_), .A2(new_n2121_), .ZN(new_n2122_));
  NAND3_X1  g1994(.A1(new_n2115_), .A2(new_n2118_), .A3(new_n2120_), .ZN(new_n2123_));
  AOI21_X1  g1995(.A(new_n2067_), .B1(new_n2122_), .B2(new_n2123_), .ZN(new_n2124_));
  INV_X1    g1996(.A(new_n2124_), .ZN(new_n2125_));
  NAND2_X1  g1997(.A1(new_n2043_), .A2(new_n2035_), .ZN(new_n2126_));
  NAND3_X1  g1998(.A1(new_n2122_), .A2(new_n2067_), .A3(new_n2123_), .ZN(new_n2127_));
  NAND3_X1  g1999(.A1(new_n2125_), .A2(new_n2126_), .A3(new_n2127_), .ZN(new_n2128_));
  NAND2_X1  g2000(.A1(G120gat), .A2(G511gat), .ZN(new_n2129_));
  INV_X1    g2001(.A(new_n2126_), .ZN(new_n2130_));
  AND3_X1   g2002(.A1(new_n2122_), .A2(new_n2067_), .A3(new_n2123_), .ZN(new_n2131_));
  OAI21_X1  g2003(.A(new_n2130_), .B1(new_n2131_), .B2(new_n2124_), .ZN(new_n2132_));
  AND3_X1   g2004(.A1(new_n2128_), .A2(new_n2129_), .A3(new_n2132_), .ZN(new_n2133_));
  AOI21_X1  g2005(.A(new_n2129_), .B1(new_n2128_), .B2(new_n2132_), .ZN(new_n2134_));
  OAI211_X1 g2006(.A(new_n2044_), .B(new_n2047_), .C1(new_n2133_), .C2(new_n2134_), .ZN(new_n2135_));
  INV_X1    g2007(.A(new_n2134_), .ZN(new_n2136_));
  NAND2_X1  g2008(.A1(new_n2047_), .A2(new_n2044_), .ZN(new_n2137_));
  NAND3_X1  g2009(.A1(new_n2128_), .A2(new_n2132_), .A3(new_n2129_), .ZN(new_n2138_));
  NAND3_X1  g2010(.A1(new_n2136_), .A2(new_n2137_), .A3(new_n2138_), .ZN(new_n2139_));
  NAND2_X1  g2011(.A1(new_n2135_), .A2(new_n2139_), .ZN(new_n2140_));
  NAND3_X1  g2012(.A1(new_n2140_), .A2(G103gat), .A3(G528gat), .ZN(new_n2141_));
  OAI211_X1 g2013(.A(new_n2135_), .B(new_n2139_), .C1(new_n243_), .C2(new_n1384_), .ZN(new_n2142_));
  NAND2_X1  g2014(.A1(new_n2057_), .A2(new_n2053_), .ZN(new_n2143_));
  AND3_X1   g2015(.A1(new_n2141_), .A2(new_n2142_), .A3(new_n2143_), .ZN(new_n2144_));
  AOI21_X1  g2016(.A(new_n2143_), .B1(new_n2141_), .B2(new_n2142_), .ZN(new_n2145_));
  NOR2_X1   g2017(.A1(new_n2144_), .A2(new_n2145_), .ZN(new_n2146_));
  XNOR2_X1  g2018(.A(new_n2066_), .B(new_n2146_), .ZN(G6200gat));
  INV_X1    g2019(.A(new_n2144_), .ZN(new_n2148_));
  AOI21_X1  g2020(.A(new_n2062_), .B1(new_n1955_), .B2(new_n2060_), .ZN(new_n2149_));
  OAI21_X1  g2021(.A(new_n2148_), .B1(new_n2149_), .B2(new_n2145_), .ZN(new_n2150_));
  NAND2_X1  g2022(.A1(G137gat), .A2(G511gat), .ZN(new_n2151_));
  NOR2_X1   g2023(.A1(new_n1084_), .A2(new_n654_), .ZN(new_n2152_));
  INV_X1    g2024(.A(new_n2152_), .ZN(new_n2153_));
  NAND2_X1  g2025(.A1(new_n2099_), .A2(new_n2098_), .ZN(new_n2154_));
  OAI21_X1  g2026(.A(new_n2069_), .B1(new_n1232_), .B2(new_n289_), .ZN(new_n2155_));
  OAI21_X1  g2027(.A(new_n2155_), .B1(new_n2076_), .B2(new_n2073_), .ZN(new_n2156_));
  OR3_X1    g2028(.A1(new_n2156_), .A2(new_n1232_), .A3(new_n363_), .ZN(new_n2157_));
  OAI21_X1  g2029(.A(new_n2156_), .B1(new_n1232_), .B2(new_n363_), .ZN(new_n2158_));
  NAND2_X1  g2030(.A1(new_n2157_), .A2(new_n2158_), .ZN(new_n2159_));
  NOR2_X1   g2031(.A1(new_n1578_), .A2(new_n443_), .ZN(new_n2160_));
  XOR2_X1   g2032(.A(new_n2159_), .B(new_n2160_), .Z(new_n2161_));
  NAND2_X1  g2033(.A1(new_n2079_), .A2(new_n2081_), .ZN(new_n2162_));
  OAI21_X1  g2034(.A(new_n2162_), .B1(new_n2082_), .B2(new_n2083_), .ZN(new_n2163_));
  XNOR2_X1  g2035(.A(new_n2161_), .B(new_n2163_), .ZN(new_n2164_));
  NOR2_X1   g2036(.A1(new_n1406_), .A2(new_n533_), .ZN(new_n2165_));
  XOR2_X1   g2037(.A(new_n2164_), .B(new_n2165_), .Z(new_n2166_));
  INV_X1    g2038(.A(new_n2166_), .ZN(new_n2167_));
  NAND3_X1  g2039(.A1(new_n2092_), .A2(KEYINPUT58), .A3(new_n2086_), .ZN(new_n2168_));
  INV_X1    g2040(.A(new_n2168_), .ZN(new_n2169_));
  AOI21_X1  g2041(.A(KEYINPUT58), .B1(new_n2092_), .B2(new_n2086_), .ZN(new_n2170_));
  OAI21_X1  g2042(.A(new_n2167_), .B1(new_n2169_), .B2(new_n2170_), .ZN(new_n2171_));
  INV_X1    g2043(.A(new_n2170_), .ZN(new_n2172_));
  NAND2_X1  g2044(.A1(new_n2172_), .A2(new_n2166_), .ZN(new_n2173_));
  NAND2_X1  g2045(.A1(new_n2171_), .A2(new_n2173_), .ZN(new_n2174_));
  OAI21_X1  g2046(.A(new_n2174_), .B1(new_n1260_), .B2(new_n648_), .ZN(new_n2175_));
  NAND4_X1  g2047(.A1(new_n2171_), .A2(G205gat), .A3(G443gat), .A4(new_n2173_), .ZN(new_n2176_));
  AOI21_X1  g2048(.A(new_n2154_), .B1(new_n2175_), .B2(new_n2176_), .ZN(new_n2177_));
  INV_X1    g2049(.A(new_n2177_), .ZN(new_n2178_));
  NAND3_X1  g2050(.A1(new_n2175_), .A2(new_n2154_), .A3(new_n2176_), .ZN(new_n2179_));
  AOI21_X1  g2051(.A(new_n2153_), .B1(new_n2178_), .B2(new_n2179_), .ZN(new_n2180_));
  INV_X1    g2052(.A(new_n2179_), .ZN(new_n2181_));
  NOR3_X1   g2053(.A1(new_n2181_), .A2(new_n2152_), .A3(new_n2177_), .ZN(new_n2182_));
  NOR2_X1   g2054(.A1(new_n2180_), .A2(new_n2182_), .ZN(new_n2183_));
  NAND2_X1  g2055(.A1(new_n2108_), .A2(new_n2105_), .ZN(new_n2184_));
  OR2_X1    g2056(.A1(new_n2183_), .A2(new_n2184_), .ZN(new_n2185_));
  NOR2_X1   g2057(.A1(new_n543_), .A2(new_n890_), .ZN(new_n2186_));
  INV_X1    g2058(.A(new_n2186_), .ZN(new_n2187_));
  NAND2_X1  g2059(.A1(new_n2183_), .A2(new_n2184_), .ZN(new_n2188_));
  AND3_X1   g2060(.A1(new_n2185_), .A2(new_n2187_), .A3(new_n2188_), .ZN(new_n2189_));
  AOI21_X1  g2061(.A(new_n2187_), .B1(new_n2185_), .B2(new_n2188_), .ZN(new_n2190_));
  AOI21_X1  g2062(.A(new_n2114_), .B1(new_n2117_), .B2(new_n2112_), .ZN(new_n2191_));
  OR3_X1    g2063(.A1(new_n2189_), .A2(new_n2190_), .A3(new_n2191_), .ZN(new_n2192_));
  NOR2_X1   g2064(.A1(new_n542_), .A2(new_n1057_), .ZN(new_n2193_));
  INV_X1    g2065(.A(new_n2193_), .ZN(new_n2194_));
  OAI21_X1  g2066(.A(new_n2191_), .B1(new_n2189_), .B2(new_n2190_), .ZN(new_n2195_));
  NAND3_X1  g2067(.A1(new_n2192_), .A2(new_n2194_), .A3(new_n2195_), .ZN(new_n2196_));
  INV_X1    g2068(.A(new_n2196_), .ZN(new_n2197_));
  AOI21_X1  g2069(.A(new_n2194_), .B1(new_n2192_), .B2(new_n2195_), .ZN(new_n2198_));
  OAI211_X1 g2070(.A(new_n2123_), .B(new_n2127_), .C1(new_n2197_), .C2(new_n2198_), .ZN(new_n2199_));
  INV_X1    g2071(.A(new_n2198_), .ZN(new_n2200_));
  NAND2_X1  g2072(.A1(new_n2127_), .A2(new_n2123_), .ZN(new_n2201_));
  NAND3_X1  g2073(.A1(new_n2200_), .A2(new_n2201_), .A3(new_n2196_), .ZN(new_n2202_));
  AOI21_X1  g2074(.A(new_n2151_), .B1(new_n2199_), .B2(new_n2202_), .ZN(new_n2203_));
  INV_X1    g2075(.A(new_n2203_), .ZN(new_n2204_));
  NAND2_X1  g2076(.A1(new_n2138_), .A2(new_n2128_), .ZN(new_n2205_));
  NAND3_X1  g2077(.A1(new_n2199_), .A2(new_n2151_), .A3(new_n2202_), .ZN(new_n2206_));
  NAND3_X1  g2078(.A1(new_n2204_), .A2(new_n2205_), .A3(new_n2206_), .ZN(new_n2207_));
  INV_X1    g2079(.A(new_n2205_), .ZN(new_n2208_));
  AND3_X1   g2080(.A1(new_n2199_), .A2(new_n2151_), .A3(new_n2202_), .ZN(new_n2209_));
  OAI21_X1  g2081(.A(new_n2208_), .B1(new_n2209_), .B2(new_n2203_), .ZN(new_n2210_));
  NOR2_X1   g2082(.A1(new_n300_), .A2(new_n1384_), .ZN(new_n2211_));
  INV_X1    g2083(.A(new_n2211_), .ZN(new_n2212_));
  NAND3_X1  g2084(.A1(new_n2207_), .A2(new_n2210_), .A3(new_n2212_), .ZN(new_n2213_));
  INV_X1    g2085(.A(new_n2213_), .ZN(new_n2214_));
  AOI21_X1  g2086(.A(new_n2212_), .B1(new_n2207_), .B2(new_n2210_), .ZN(new_n2215_));
  OAI211_X1 g2087(.A(new_n2139_), .B(new_n2142_), .C1(new_n2214_), .C2(new_n2215_), .ZN(new_n2216_));
  INV_X1    g2088(.A(new_n2215_), .ZN(new_n2217_));
  NAND2_X1  g2089(.A1(new_n2142_), .A2(new_n2139_), .ZN(new_n2218_));
  NAND3_X1  g2090(.A1(new_n2217_), .A2(new_n2218_), .A3(new_n2213_), .ZN(new_n2219_));
  AND2_X1   g2091(.A1(new_n2216_), .A2(new_n2219_), .ZN(new_n2220_));
  XNOR2_X1  g2092(.A(new_n2150_), .B(new_n2220_), .ZN(G6210gat));
  AOI21_X1  g2093(.A(new_n2144_), .B1(new_n2066_), .B2(new_n2146_), .ZN(new_n2222_));
  INV_X1    g2094(.A(new_n2216_), .ZN(new_n2223_));
  OAI21_X1  g2095(.A(new_n2219_), .B1(new_n2222_), .B2(new_n2223_), .ZN(new_n2224_));
  NOR2_X1   g2096(.A1(new_n2183_), .A2(new_n2184_), .ZN(new_n2225_));
  OAI21_X1  g2097(.A(new_n2188_), .B1(new_n2225_), .B2(new_n2186_), .ZN(new_n2226_));
  INV_X1    g2098(.A(new_n2226_), .ZN(new_n2227_));
  NAND2_X1  g2099(.A1(new_n2092_), .A2(new_n2086_), .ZN(new_n2228_));
  NAND2_X1  g2100(.A1(new_n2166_), .A2(new_n2228_), .ZN(new_n2229_));
  AND2_X1   g2101(.A1(new_n2175_), .A2(new_n2229_), .ZN(new_n2230_));
  OR2_X1    g2102(.A1(new_n2164_), .A2(new_n2165_), .ZN(new_n2231_));
  NAND2_X1  g2103(.A1(new_n2161_), .A2(new_n2163_), .ZN(new_n2232_));
  NAND2_X1  g2104(.A1(new_n2231_), .A2(new_n2232_), .ZN(new_n2233_));
  OAI21_X1  g2105(.A(new_n2158_), .B1(new_n2159_), .B2(new_n2160_), .ZN(new_n2234_));
  OR3_X1    g2106(.A1(new_n2234_), .A2(new_n1232_), .A3(new_n443_), .ZN(new_n2235_));
  OAI21_X1  g2107(.A(new_n2234_), .B1(new_n1232_), .B2(new_n443_), .ZN(new_n2236_));
  NAND2_X1  g2108(.A1(new_n2235_), .A2(new_n2236_), .ZN(new_n2237_));
  NOR2_X1   g2109(.A1(new_n1578_), .A2(new_n533_), .ZN(new_n2238_));
  OR2_X1    g2110(.A1(new_n2237_), .A2(new_n2238_), .ZN(new_n2239_));
  NAND2_X1  g2111(.A1(new_n2237_), .A2(new_n2238_), .ZN(new_n2240_));
  NAND2_X1  g2112(.A1(new_n2239_), .A2(new_n2240_), .ZN(new_n2241_));
  XOR2_X1   g2113(.A(new_n2233_), .B(new_n2241_), .Z(new_n2242_));
  NOR2_X1   g2114(.A1(new_n1406_), .A2(new_n648_), .ZN(new_n2243_));
  XNOR2_X1  g2115(.A(new_n2242_), .B(new_n2243_), .ZN(new_n2244_));
  NOR2_X1   g2116(.A1(new_n2230_), .A2(new_n2244_), .ZN(new_n2245_));
  INV_X1    g2117(.A(new_n2245_), .ZN(new_n2246_));
  NAND2_X1  g2118(.A1(new_n2230_), .A2(new_n2244_), .ZN(new_n2247_));
  OAI211_X1 g2119(.A(new_n2246_), .B(new_n2247_), .C1(new_n1260_), .C2(new_n654_), .ZN(new_n2248_));
  AND2_X1   g2120(.A1(new_n2230_), .A2(new_n2244_), .ZN(new_n2249_));
  OAI211_X1 g2121(.A(G205gat), .B(G460gat), .C1(new_n2249_), .C2(new_n2245_), .ZN(new_n2250_));
  NAND2_X1  g2122(.A1(new_n2248_), .A2(new_n2250_), .ZN(new_n2251_));
  INV_X1    g2123(.A(new_n2182_), .ZN(new_n2252_));
  NAND3_X1  g2124(.A1(new_n2251_), .A2(new_n2179_), .A3(new_n2252_), .ZN(new_n2253_));
  NOR2_X1   g2125(.A1(new_n1084_), .A2(new_n890_), .ZN(new_n2254_));
  INV_X1    g2126(.A(new_n2254_), .ZN(new_n2255_));
  OAI211_X1 g2127(.A(new_n2248_), .B(new_n2250_), .C1(new_n2181_), .C2(new_n2182_), .ZN(new_n2256_));
  NAND3_X1  g2128(.A1(new_n2253_), .A2(new_n2255_), .A3(new_n2256_), .ZN(new_n2257_));
  INV_X1    g2129(.A(new_n2257_), .ZN(new_n2258_));
  AOI21_X1  g2130(.A(new_n2255_), .B1(new_n2253_), .B2(new_n2256_), .ZN(new_n2259_));
  OAI21_X1  g2131(.A(new_n2227_), .B1(new_n2258_), .B2(new_n2259_), .ZN(new_n2260_));
  INV_X1    g2132(.A(new_n2259_), .ZN(new_n2261_));
  NAND3_X1  g2133(.A1(new_n2261_), .A2(new_n2226_), .A3(new_n2257_), .ZN(new_n2262_));
  NAND2_X1  g2134(.A1(new_n2260_), .A2(new_n2262_), .ZN(new_n2263_));
  NOR2_X1   g2135(.A1(new_n543_), .A2(new_n1057_), .ZN(new_n2264_));
  NAND2_X1  g2136(.A1(new_n2263_), .A2(new_n2264_), .ZN(new_n2265_));
  OAI211_X1 g2137(.A(new_n2260_), .B(new_n2262_), .C1(new_n543_), .C2(new_n1057_), .ZN(new_n2266_));
  NAND2_X1  g2138(.A1(new_n2265_), .A2(new_n2266_), .ZN(new_n2267_));
  NAND3_X1  g2139(.A1(new_n2267_), .A2(new_n2192_), .A3(new_n2196_), .ZN(new_n2268_));
  NOR2_X1   g2140(.A1(new_n542_), .A2(new_n1218_), .ZN(new_n2269_));
  INV_X1    g2141(.A(new_n2269_), .ZN(new_n2270_));
  NAND2_X1  g2142(.A1(new_n2196_), .A2(new_n2192_), .ZN(new_n2271_));
  NAND3_X1  g2143(.A1(new_n2265_), .A2(new_n2271_), .A3(new_n2266_), .ZN(new_n2272_));
  NAND3_X1  g2144(.A1(new_n2268_), .A2(new_n2270_), .A3(new_n2272_), .ZN(new_n2273_));
  INV_X1    g2145(.A(new_n2273_), .ZN(new_n2274_));
  AOI21_X1  g2146(.A(new_n2270_), .B1(new_n2268_), .B2(new_n2272_), .ZN(new_n2275_));
  NOR2_X1   g2147(.A1(new_n2274_), .A2(new_n2275_), .ZN(new_n2276_));
  NAND2_X1  g2148(.A1(new_n2206_), .A2(new_n2202_), .ZN(new_n2277_));
  NAND2_X1  g2149(.A1(new_n2276_), .A2(new_n2277_), .ZN(new_n2278_));
  NOR2_X1   g2150(.A1(new_n377_), .A2(new_n1384_), .ZN(new_n2279_));
  INV_X1    g2151(.A(new_n2279_), .ZN(new_n2280_));
  OAI211_X1 g2152(.A(new_n2202_), .B(new_n2206_), .C1(new_n2274_), .C2(new_n2275_), .ZN(new_n2281_));
  NAND3_X1  g2153(.A1(new_n2278_), .A2(new_n2280_), .A3(new_n2281_), .ZN(new_n2282_));
  INV_X1    g2154(.A(new_n2282_), .ZN(new_n2283_));
  AOI21_X1  g2155(.A(new_n2280_), .B1(new_n2278_), .B2(new_n2281_), .ZN(new_n2284_));
  NOR2_X1   g2156(.A1(new_n2283_), .A2(new_n2284_), .ZN(new_n2285_));
  NAND2_X1  g2157(.A1(new_n2213_), .A2(new_n2207_), .ZN(new_n2286_));
  NAND2_X1  g2158(.A1(new_n2285_), .A2(new_n2286_), .ZN(new_n2287_));
  OAI211_X1 g2159(.A(new_n2207_), .B(new_n2213_), .C1(new_n2283_), .C2(new_n2284_), .ZN(new_n2288_));
  AND2_X1   g2160(.A1(new_n2287_), .A2(new_n2288_), .ZN(new_n2289_));
  XNOR2_X1  g2161(.A(new_n2224_), .B(new_n2289_), .ZN(G6220gat));
  INV_X1    g2162(.A(new_n2219_), .ZN(new_n2291_));
  AOI21_X1  g2163(.A(new_n2291_), .B1(new_n2150_), .B2(new_n2220_), .ZN(new_n2292_));
  INV_X1    g2164(.A(new_n2288_), .ZN(new_n2293_));
  OAI21_X1  g2165(.A(new_n2287_), .B1(new_n2292_), .B2(new_n2293_), .ZN(new_n2294_));
  NOR2_X1   g2166(.A1(new_n542_), .A2(new_n1384_), .ZN(new_n2295_));
  INV_X1    g2167(.A(KEYINPUT60), .ZN(new_n2296_));
  NAND2_X1  g2168(.A1(new_n2248_), .A2(new_n2246_), .ZN(new_n2297_));
  OR2_X1    g2169(.A1(new_n2242_), .A2(new_n2243_), .ZN(new_n2298_));
  NAND3_X1  g2170(.A1(new_n2233_), .A2(new_n2239_), .A3(new_n2240_), .ZN(new_n2299_));
  NAND2_X1  g2171(.A1(new_n2298_), .A2(new_n2299_), .ZN(new_n2300_));
  NAND2_X1  g2172(.A1(new_n2239_), .A2(new_n2236_), .ZN(new_n2301_));
  NAND2_X1  g2173(.A1(G256gat), .A2(G426gat), .ZN(new_n2302_));
  OR2_X1    g2174(.A1(new_n2301_), .A2(new_n2302_), .ZN(new_n2303_));
  NAND2_X1  g2175(.A1(new_n2301_), .A2(new_n2302_), .ZN(new_n2304_));
  NAND2_X1  g2176(.A1(new_n2303_), .A2(new_n2304_), .ZN(new_n2305_));
  NOR2_X1   g2177(.A1(new_n1578_), .A2(new_n648_), .ZN(new_n2306_));
  OR2_X1    g2178(.A1(new_n2305_), .A2(new_n2306_), .ZN(new_n2307_));
  NAND2_X1  g2179(.A1(new_n2305_), .A2(new_n2306_), .ZN(new_n2308_));
  NAND3_X1  g2180(.A1(new_n2300_), .A2(new_n2307_), .A3(new_n2308_), .ZN(new_n2309_));
  NAND2_X1  g2181(.A1(new_n2307_), .A2(new_n2308_), .ZN(new_n2310_));
  NAND3_X1  g2182(.A1(new_n2298_), .A2(new_n2299_), .A3(new_n2310_), .ZN(new_n2311_));
  OAI211_X1 g2183(.A(new_n2309_), .B(new_n2311_), .C1(new_n1406_), .C2(new_n654_), .ZN(new_n2312_));
  NAND2_X1  g2184(.A1(new_n2309_), .A2(new_n2311_), .ZN(new_n2313_));
  NAND3_X1  g2185(.A1(new_n2313_), .A2(G222gat), .A3(G460gat), .ZN(new_n2314_));
  NAND3_X1  g2186(.A1(new_n2297_), .A2(new_n2312_), .A3(new_n2314_), .ZN(new_n2315_));
  NAND2_X1  g2187(.A1(G205gat), .A2(G477gat), .ZN(new_n2316_));
  XNOR2_X1  g2188(.A(new_n2316_), .B(KEYINPUT59), .ZN(new_n2317_));
  INV_X1    g2189(.A(new_n2317_), .ZN(new_n2318_));
  NAND2_X1  g2190(.A1(new_n2314_), .A2(new_n2312_), .ZN(new_n2319_));
  NAND3_X1  g2191(.A1(new_n2319_), .A2(new_n2248_), .A3(new_n2246_), .ZN(new_n2320_));
  NAND3_X1  g2192(.A1(new_n2315_), .A2(new_n2318_), .A3(new_n2320_), .ZN(new_n2321_));
  INV_X1    g2193(.A(new_n2321_), .ZN(new_n2322_));
  AOI21_X1  g2194(.A(new_n2318_), .B1(new_n2315_), .B2(new_n2320_), .ZN(new_n2323_));
  OAI21_X1  g2195(.A(new_n2296_), .B1(new_n2322_), .B2(new_n2323_), .ZN(new_n2324_));
  INV_X1    g2196(.A(new_n2323_), .ZN(new_n2325_));
  NAND3_X1  g2197(.A1(new_n2325_), .A2(KEYINPUT60), .A3(new_n2321_), .ZN(new_n2326_));
  NAND2_X1  g2198(.A1(new_n2257_), .A2(new_n2256_), .ZN(new_n2327_));
  NAND3_X1  g2199(.A1(new_n2324_), .A2(new_n2326_), .A3(new_n2327_), .ZN(new_n2328_));
  NAND2_X1  g2200(.A1(G188gat), .A2(G494gat), .ZN(new_n2329_));
  OAI211_X1 g2201(.A(new_n2256_), .B(new_n2257_), .C1(new_n2322_), .C2(new_n2323_), .ZN(new_n2330_));
  NAND3_X1  g2202(.A1(new_n2328_), .A2(new_n2329_), .A3(new_n2330_), .ZN(new_n2331_));
  INV_X1    g2203(.A(new_n2331_), .ZN(new_n2332_));
  AND2_X1   g2204(.A1(new_n2266_), .A2(new_n2262_), .ZN(new_n2333_));
  AOI21_X1  g2205(.A(new_n2329_), .B1(new_n2328_), .B2(new_n2330_), .ZN(new_n2334_));
  OR3_X1    g2206(.A1(new_n2332_), .A2(new_n2333_), .A3(new_n2334_), .ZN(new_n2335_));
  NOR2_X1   g2207(.A1(new_n543_), .A2(new_n1218_), .ZN(new_n2336_));
  INV_X1    g2208(.A(new_n2336_), .ZN(new_n2337_));
  OAI21_X1  g2209(.A(new_n2333_), .B1(new_n2332_), .B2(new_n2334_), .ZN(new_n2338_));
  NAND3_X1  g2210(.A1(new_n2335_), .A2(new_n2337_), .A3(new_n2338_), .ZN(new_n2339_));
  INV_X1    g2211(.A(new_n2339_), .ZN(new_n2340_));
  AOI21_X1  g2212(.A(new_n2337_), .B1(new_n2335_), .B2(new_n2338_), .ZN(new_n2341_));
  NOR2_X1   g2213(.A1(new_n2340_), .A2(new_n2341_), .ZN(new_n2342_));
  NAND2_X1  g2214(.A1(new_n2273_), .A2(new_n2272_), .ZN(new_n2343_));
  NOR2_X1   g2215(.A1(new_n2342_), .A2(new_n2343_), .ZN(new_n2344_));
  INV_X1    g2216(.A(new_n2341_), .ZN(new_n2345_));
  NAND2_X1  g2217(.A1(new_n2345_), .A2(new_n2339_), .ZN(new_n2346_));
  INV_X1    g2218(.A(new_n2343_), .ZN(new_n2347_));
  NOR2_X1   g2219(.A1(new_n2346_), .A2(new_n2347_), .ZN(new_n2348_));
  OAI21_X1  g2220(.A(new_n2295_), .B1(new_n2344_), .B2(new_n2348_), .ZN(new_n2349_));
  NAND2_X1  g2221(.A1(new_n2342_), .A2(new_n2343_), .ZN(new_n2350_));
  NAND2_X1  g2222(.A1(new_n2346_), .A2(new_n2347_), .ZN(new_n2351_));
  INV_X1    g2223(.A(new_n2295_), .ZN(new_n2352_));
  NAND3_X1  g2224(.A1(new_n2350_), .A2(new_n2351_), .A3(new_n2352_), .ZN(new_n2353_));
  NAND2_X1  g2225(.A1(new_n2349_), .A2(new_n2353_), .ZN(new_n2354_));
  NAND2_X1  g2226(.A1(new_n2282_), .A2(new_n2278_), .ZN(new_n2355_));
  XNOR2_X1  g2227(.A(new_n2354_), .B(new_n2355_), .ZN(new_n2356_));
  XNOR2_X1  g2228(.A(new_n2294_), .B(new_n2356_), .ZN(G6230gat));
  INV_X1    g2229(.A(new_n2354_), .ZN(new_n2358_));
  NAND2_X1  g2230(.A1(new_n2358_), .A2(new_n2355_), .ZN(new_n2359_));
  INV_X1    g2231(.A(new_n2359_), .ZN(new_n2360_));
  AOI21_X1  g2232(.A(new_n2360_), .B1(new_n2294_), .B2(new_n2356_), .ZN(new_n2361_));
  AND2_X1   g2233(.A1(new_n2331_), .A2(new_n2328_), .ZN(new_n2362_));
  NAND2_X1  g2234(.A1(new_n2312_), .A2(new_n2309_), .ZN(new_n2363_));
  INV_X1    g2235(.A(KEYINPUT61), .ZN(new_n2364_));
  NAND2_X1  g2236(.A1(new_n2363_), .A2(new_n2364_), .ZN(new_n2365_));
  NAND3_X1  g2237(.A1(new_n2312_), .A2(KEYINPUT61), .A3(new_n2309_), .ZN(new_n2366_));
  NAND2_X1  g2238(.A1(new_n2307_), .A2(new_n2304_), .ZN(new_n2367_));
  OAI21_X1  g2239(.A(new_n2367_), .B1(new_n1232_), .B2(new_n648_), .ZN(new_n2368_));
  NAND4_X1  g2240(.A1(new_n2307_), .A2(G256gat), .A3(G443gat), .A4(new_n2304_), .ZN(new_n2369_));
  NAND2_X1  g2241(.A1(new_n2368_), .A2(new_n2369_), .ZN(new_n2370_));
  NOR2_X1   g2242(.A1(new_n1578_), .A2(new_n654_), .ZN(new_n2371_));
  XOR2_X1   g2243(.A(new_n2370_), .B(new_n2371_), .Z(new_n2372_));
  NAND3_X1  g2244(.A1(new_n2365_), .A2(new_n2366_), .A3(new_n2372_), .ZN(new_n2373_));
  INV_X1    g2245(.A(new_n2373_), .ZN(new_n2374_));
  NOR2_X1   g2246(.A1(new_n1406_), .A2(new_n890_), .ZN(new_n2375_));
  AOI21_X1  g2247(.A(new_n2372_), .B1(new_n2365_), .B2(new_n2366_), .ZN(new_n2376_));
  OR3_X1    g2248(.A1(new_n2374_), .A2(new_n2375_), .A3(new_n2376_), .ZN(new_n2377_));
  OAI21_X1  g2249(.A(new_n2375_), .B1(new_n2374_), .B2(new_n2376_), .ZN(new_n2378_));
  NAND2_X1  g2250(.A1(new_n2377_), .A2(new_n2378_), .ZN(new_n2379_));
  AND2_X1   g2251(.A1(new_n2321_), .A2(new_n2315_), .ZN(new_n2380_));
  OR2_X1    g2252(.A1(new_n2379_), .A2(new_n2380_), .ZN(new_n2381_));
  NAND2_X1  g2253(.A1(G205gat), .A2(G494gat), .ZN(new_n2382_));
  NAND2_X1  g2254(.A1(new_n2379_), .A2(new_n2380_), .ZN(new_n2383_));
  NAND3_X1  g2255(.A1(new_n2381_), .A2(new_n2382_), .A3(new_n2383_), .ZN(new_n2384_));
  INV_X1    g2256(.A(new_n2384_), .ZN(new_n2385_));
  AOI21_X1  g2257(.A(new_n2382_), .B1(new_n2381_), .B2(new_n2383_), .ZN(new_n2386_));
  OR3_X1    g2258(.A1(new_n2362_), .A2(new_n2385_), .A3(new_n2386_), .ZN(new_n2387_));
  NAND2_X1  g2259(.A1(G188gat), .A2(G511gat), .ZN(new_n2388_));
  OAI21_X1  g2260(.A(new_n2362_), .B1(new_n2385_), .B2(new_n2386_), .ZN(new_n2389_));
  NAND3_X1  g2261(.A1(new_n2387_), .A2(new_n2388_), .A3(new_n2389_), .ZN(new_n2390_));
  INV_X1    g2262(.A(new_n2390_), .ZN(new_n2391_));
  AOI21_X1  g2263(.A(new_n2388_), .B1(new_n2387_), .B2(new_n2389_), .ZN(new_n2392_));
  NOR2_X1   g2264(.A1(new_n2391_), .A2(new_n2392_), .ZN(new_n2393_));
  NAND2_X1  g2265(.A1(new_n2339_), .A2(new_n2335_), .ZN(new_n2394_));
  OR2_X1    g2266(.A1(new_n2393_), .A2(new_n2394_), .ZN(new_n2395_));
  NAND2_X1  g2267(.A1(new_n2393_), .A2(new_n2394_), .ZN(new_n2396_));
  NAND2_X1  g2268(.A1(new_n2395_), .A2(new_n2396_), .ZN(new_n2397_));
  NAND3_X1  g2269(.A1(new_n2397_), .A2(G171gat), .A3(G528gat), .ZN(new_n2398_));
  OAI211_X1 g2270(.A(new_n2395_), .B(new_n2396_), .C1(new_n543_), .C2(new_n1384_), .ZN(new_n2399_));
  NAND2_X1  g2271(.A1(new_n2398_), .A2(new_n2399_), .ZN(new_n2400_));
  NAND3_X1  g2272(.A1(new_n2400_), .A2(new_n2350_), .A3(new_n2353_), .ZN(new_n2401_));
  NAND2_X1  g2273(.A1(new_n2353_), .A2(new_n2350_), .ZN(new_n2402_));
  NAND3_X1  g2274(.A1(new_n2398_), .A2(new_n2399_), .A3(new_n2402_), .ZN(new_n2403_));
  NAND2_X1  g2275(.A1(new_n2401_), .A2(new_n2403_), .ZN(new_n2404_));
  XNOR2_X1  g2276(.A(new_n2361_), .B(new_n2404_), .ZN(G6240gat));
  INV_X1    g2277(.A(new_n2403_), .ZN(new_n2406_));
  INV_X1    g2278(.A(new_n2287_), .ZN(new_n2407_));
  AOI21_X1  g2279(.A(new_n2407_), .B1(new_n2224_), .B2(new_n2289_), .ZN(new_n2408_));
  NOR2_X1   g2280(.A1(new_n2358_), .A2(new_n2355_), .ZN(new_n2409_));
  OAI21_X1  g2281(.A(new_n2359_), .B1(new_n2408_), .B2(new_n2409_), .ZN(new_n2410_));
  AOI21_X1  g2282(.A(new_n2406_), .B1(new_n2410_), .B2(new_n2401_), .ZN(new_n2411_));
  NAND2_X1  g2283(.A1(new_n2377_), .A2(new_n2373_), .ZN(new_n2412_));
  OAI21_X1  g2284(.A(new_n2368_), .B1(new_n2370_), .B2(new_n2371_), .ZN(new_n2413_));
  OR3_X1    g2285(.A1(new_n2413_), .A2(new_n1232_), .A3(new_n654_), .ZN(new_n2414_));
  OAI21_X1  g2286(.A(new_n2413_), .B1(new_n1232_), .B2(new_n654_), .ZN(new_n2415_));
  NAND2_X1  g2287(.A1(new_n2414_), .A2(new_n2415_), .ZN(new_n2416_));
  NOR2_X1   g2288(.A1(new_n1578_), .A2(new_n890_), .ZN(new_n2417_));
  XOR2_X1   g2289(.A(new_n2416_), .B(new_n2417_), .Z(new_n2418_));
  XNOR2_X1  g2290(.A(new_n2412_), .B(new_n2418_), .ZN(new_n2419_));
  NOR2_X1   g2291(.A1(new_n1406_), .A2(new_n1057_), .ZN(new_n2420_));
  XNOR2_X1  g2292(.A(new_n2419_), .B(new_n2420_), .ZN(new_n2421_));
  AND2_X1   g2293(.A1(new_n2384_), .A2(new_n2381_), .ZN(new_n2422_));
  XNOR2_X1  g2294(.A(new_n2421_), .B(new_n2422_), .ZN(new_n2423_));
  NOR2_X1   g2295(.A1(new_n1260_), .A2(new_n1218_), .ZN(new_n2424_));
  XNOR2_X1  g2296(.A(new_n2423_), .B(new_n2424_), .ZN(new_n2425_));
  NAND2_X1  g2297(.A1(new_n2390_), .A2(new_n2387_), .ZN(new_n2426_));
  XNOR2_X1  g2298(.A(new_n2425_), .B(new_n2426_), .ZN(new_n2427_));
  INV_X1    g2299(.A(new_n2427_), .ZN(new_n2428_));
  NAND3_X1  g2300(.A1(new_n2428_), .A2(G188gat), .A3(G528gat), .ZN(new_n2429_));
  OAI21_X1  g2301(.A(new_n2427_), .B1(new_n1084_), .B2(new_n1384_), .ZN(new_n2430_));
  NAND2_X1  g2302(.A1(new_n2429_), .A2(new_n2430_), .ZN(new_n2431_));
  NAND2_X1  g2303(.A1(new_n2399_), .A2(new_n2396_), .ZN(new_n2432_));
  INV_X1    g2304(.A(new_n2432_), .ZN(new_n2433_));
  XNOR2_X1  g2305(.A(new_n2431_), .B(new_n2433_), .ZN(new_n2434_));
  NAND2_X1  g2306(.A1(new_n2411_), .A2(new_n2434_), .ZN(new_n2435_));
  OAI21_X1  g2307(.A(new_n2403_), .B1(new_n2361_), .B2(new_n2404_), .ZN(new_n2436_));
  XNOR2_X1  g2308(.A(new_n2431_), .B(new_n2432_), .ZN(new_n2437_));
  NAND2_X1  g2309(.A1(new_n2436_), .A2(new_n2437_), .ZN(new_n2438_));
  NAND2_X1  g2310(.A1(new_n2435_), .A2(new_n2438_), .ZN(G6250gat));
  INV_X1    g2311(.A(new_n2431_), .ZN(new_n2440_));
  NAND2_X1  g2312(.A1(new_n2440_), .A2(new_n2432_), .ZN(new_n2441_));
  NAND2_X1  g2313(.A1(new_n2438_), .A2(new_n2441_), .ZN(new_n2442_));
  NAND3_X1  g2314(.A1(new_n2440_), .A2(KEYINPUT62), .A3(new_n2432_), .ZN(new_n2443_));
  INV_X1    g2315(.A(KEYINPUT62), .ZN(new_n2444_));
  OAI21_X1  g2316(.A(new_n2444_), .B1(new_n2431_), .B2(new_n2433_), .ZN(new_n2445_));
  NAND2_X1  g2317(.A1(new_n2443_), .A2(new_n2445_), .ZN(new_n2446_));
  AND2_X1   g2318(.A1(new_n2438_), .A2(new_n2446_), .ZN(new_n2447_));
  INV_X1    g2319(.A(new_n2426_), .ZN(new_n2448_));
  OAI21_X1  g2320(.A(new_n2430_), .B1(new_n2448_), .B2(new_n2425_), .ZN(new_n2449_));
  NOR2_X1   g2321(.A1(new_n2423_), .A2(new_n2424_), .ZN(new_n2450_));
  NOR2_X1   g2322(.A1(new_n2421_), .A2(new_n2422_), .ZN(new_n2451_));
  NOR2_X1   g2323(.A1(new_n2450_), .A2(new_n2451_), .ZN(new_n2452_));
  NAND2_X1  g2324(.A1(new_n2412_), .A2(new_n2418_), .ZN(new_n2453_));
  OAI21_X1  g2325(.A(new_n2453_), .B1(new_n2419_), .B2(new_n2420_), .ZN(new_n2454_));
  OAI21_X1  g2326(.A(new_n2415_), .B1(new_n2416_), .B2(new_n2417_), .ZN(new_n2455_));
  OR3_X1    g2327(.A1(new_n2455_), .A2(new_n1232_), .A3(new_n890_), .ZN(new_n2456_));
  OAI21_X1  g2328(.A(new_n2455_), .B1(new_n1232_), .B2(new_n890_), .ZN(new_n2457_));
  NAND2_X1  g2329(.A1(new_n2456_), .A2(new_n2457_), .ZN(new_n2458_));
  NOR2_X1   g2330(.A1(new_n1578_), .A2(new_n1057_), .ZN(new_n2459_));
  XNOR2_X1  g2331(.A(new_n2458_), .B(new_n2459_), .ZN(new_n2460_));
  XOR2_X1   g2332(.A(new_n2454_), .B(new_n2460_), .Z(new_n2461_));
  NOR2_X1   g2333(.A1(new_n1406_), .A2(new_n1218_), .ZN(new_n2462_));
  XNOR2_X1  g2334(.A(new_n2461_), .B(new_n2462_), .ZN(new_n2463_));
  OR2_X1    g2335(.A1(new_n2452_), .A2(new_n2463_), .ZN(new_n2464_));
  NAND2_X1  g2336(.A1(new_n2452_), .A2(new_n2463_), .ZN(new_n2465_));
  NAND2_X1  g2337(.A1(new_n2464_), .A2(new_n2465_), .ZN(new_n2466_));
  NAND2_X1  g2338(.A1(G205gat), .A2(G528gat), .ZN(new_n2467_));
  XNOR2_X1  g2339(.A(new_n2466_), .B(new_n2467_), .ZN(new_n2468_));
  NOR2_X1   g2340(.A1(new_n2449_), .A2(new_n2468_), .ZN(new_n2469_));
  INV_X1    g2341(.A(new_n2469_), .ZN(new_n2470_));
  NAND2_X1  g2342(.A1(new_n2449_), .A2(new_n2468_), .ZN(new_n2471_));
  NAND2_X1  g2343(.A1(new_n2470_), .A2(new_n2471_), .ZN(new_n2472_));
  MUX2_X1   g2344(.A(new_n2442_), .B(new_n2447_), .S(new_n2472_), .Z(G6260gat));
  OAI211_X1 g2345(.A(new_n2471_), .B(new_n2446_), .C1(new_n2411_), .C2(new_n2434_), .ZN(new_n2474_));
  NAND2_X1  g2346(.A1(new_n2474_), .A2(new_n2470_), .ZN(new_n2475_));
  OR2_X1    g2347(.A1(new_n2461_), .A2(new_n2462_), .ZN(new_n2476_));
  INV_X1    g2348(.A(new_n2454_), .ZN(new_n2477_));
  OR2_X1    g2349(.A1(new_n2477_), .A2(new_n2460_), .ZN(new_n2478_));
  NAND2_X1  g2350(.A1(new_n2476_), .A2(new_n2478_), .ZN(new_n2479_));
  OAI21_X1  g2351(.A(new_n2457_), .B1(new_n2458_), .B2(new_n2459_), .ZN(new_n2480_));
  NAND2_X1  g2352(.A1(G256gat), .A2(G494gat), .ZN(new_n2481_));
  XNOR2_X1  g2353(.A(new_n2480_), .B(new_n2481_), .ZN(new_n2482_));
  NOR2_X1   g2354(.A1(new_n1578_), .A2(new_n1218_), .ZN(new_n2483_));
  XOR2_X1   g2355(.A(new_n2482_), .B(new_n2483_), .Z(new_n2484_));
  XNOR2_X1  g2356(.A(new_n2479_), .B(new_n2484_), .ZN(new_n2485_));
  NOR2_X1   g2357(.A1(new_n1406_), .A2(new_n1384_), .ZN(new_n2486_));
  XOR2_X1   g2358(.A(new_n2485_), .B(new_n2486_), .Z(new_n2487_));
  NAND3_X1  g2359(.A1(new_n2464_), .A2(new_n2467_), .A3(new_n2465_), .ZN(new_n2488_));
  NAND2_X1  g2360(.A1(new_n2488_), .A2(new_n2464_), .ZN(new_n2489_));
  OR2_X1    g2361(.A1(new_n2487_), .A2(new_n2489_), .ZN(new_n2490_));
  NAND2_X1  g2362(.A1(new_n2487_), .A2(new_n2489_), .ZN(new_n2491_));
  AND2_X1   g2363(.A1(new_n2490_), .A2(new_n2491_), .ZN(new_n2492_));
  XOR2_X1   g2364(.A(new_n2475_), .B(new_n2492_), .Z(G6270gat));
  NAND3_X1  g2365(.A1(new_n2474_), .A2(new_n2470_), .A3(new_n2492_), .ZN(new_n2494_));
  NAND2_X1  g2366(.A1(new_n2479_), .A2(new_n2484_), .ZN(new_n2495_));
  OAI21_X1  g2367(.A(new_n2495_), .B1(new_n2485_), .B2(new_n2486_), .ZN(new_n2496_));
  OR2_X1    g2368(.A1(new_n2482_), .A2(new_n2483_), .ZN(new_n2497_));
  NAND2_X1  g2369(.A1(new_n2480_), .A2(new_n2481_), .ZN(new_n2498_));
  NAND2_X1  g2370(.A1(new_n2497_), .A2(new_n2498_), .ZN(new_n2499_));
  OAI21_X1  g2371(.A(new_n2499_), .B1(new_n1232_), .B2(new_n1218_), .ZN(new_n2500_));
  NAND4_X1  g2372(.A1(new_n2497_), .A2(G256gat), .A3(G511gat), .A4(new_n2498_), .ZN(new_n2501_));
  NAND2_X1  g2373(.A1(new_n2500_), .A2(new_n2501_), .ZN(new_n2502_));
  NAND2_X1  g2374(.A1(G239gat), .A2(G528gat), .ZN(new_n2503_));
  XNOR2_X1  g2375(.A(new_n2502_), .B(new_n2503_), .ZN(new_n2504_));
  OR2_X1    g2376(.A1(new_n2496_), .A2(new_n2504_), .ZN(new_n2505_));
  NAND2_X1  g2377(.A1(new_n2496_), .A2(new_n2504_), .ZN(new_n2506_));
  NAND2_X1  g2378(.A1(new_n2505_), .A2(new_n2506_), .ZN(new_n2507_));
  NAND3_X1  g2379(.A1(new_n2494_), .A2(new_n2491_), .A3(new_n2507_), .ZN(new_n2508_));
  INV_X1    g2380(.A(new_n2441_), .ZN(new_n2509_));
  AOI21_X1  g2381(.A(new_n2509_), .B1(new_n2436_), .B2(new_n2437_), .ZN(new_n2510_));
  OAI211_X1 g2382(.A(new_n2471_), .B(new_n2491_), .C1(new_n2510_), .C2(new_n2469_), .ZN(new_n2511_));
  AND3_X1   g2383(.A1(new_n2490_), .A2(new_n2506_), .A3(new_n2505_), .ZN(new_n2512_));
  NAND2_X1  g2384(.A1(new_n2511_), .A2(new_n2512_), .ZN(new_n2513_));
  NAND2_X1  g2385(.A1(new_n2508_), .A2(new_n2513_), .ZN(new_n2514_));
  NAND2_X1  g2386(.A1(new_n2514_), .A2(KEYINPUT63), .ZN(new_n2515_));
  INV_X1    g2387(.A(KEYINPUT63), .ZN(new_n2516_));
  NAND3_X1  g2388(.A1(new_n2508_), .A2(new_n2516_), .A3(new_n2513_), .ZN(new_n2517_));
  NAND2_X1  g2389(.A1(new_n2515_), .A2(new_n2517_), .ZN(G6280gat));
  NAND3_X1  g2390(.A1(new_n2500_), .A2(new_n2501_), .A3(new_n2503_), .ZN(new_n2519_));
  NAND2_X1  g2391(.A1(new_n2519_), .A2(new_n2500_), .ZN(new_n2520_));
  INV_X1    g2392(.A(new_n2520_), .ZN(new_n2521_));
  NOR2_X1   g2393(.A1(new_n1232_), .A2(new_n1384_), .ZN(new_n2522_));
  NOR2_X1   g2394(.A1(new_n2521_), .A2(new_n2522_), .ZN(new_n2523_));
  NAND2_X1  g2395(.A1(new_n2513_), .A2(new_n2506_), .ZN(new_n2524_));
  NAND2_X1  g2396(.A1(new_n2521_), .A2(new_n2522_), .ZN(new_n2525_));
  AOI21_X1  g2397(.A(new_n2523_), .B1(new_n2524_), .B2(new_n2525_), .ZN(G6287gat));
  INV_X1    g2398(.A(new_n2525_), .ZN(new_n2527_));
  NOR2_X1   g2399(.A1(new_n2527_), .A2(new_n2523_), .ZN(new_n2528_));
  AOI21_X1  g2400(.A(new_n2528_), .B1(new_n2513_), .B2(new_n2506_), .ZN(new_n2529_));
  INV_X1    g2401(.A(new_n2506_), .ZN(new_n2530_));
  NAND2_X1  g2402(.A1(new_n2494_), .A2(new_n2491_), .ZN(new_n2531_));
  AOI21_X1  g2403(.A(new_n2530_), .B1(new_n2531_), .B2(new_n2505_), .ZN(new_n2532_));
  AOI21_X1  g2404(.A(new_n2529_), .B1(new_n2528_), .B2(new_n2532_), .ZN(G6288gat));
endmodule


