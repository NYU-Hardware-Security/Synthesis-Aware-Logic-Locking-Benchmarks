//Secret key is'1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_c2670" written by ABC on Wed Oct 26 13:56:14 2022

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6,
    G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26,
    G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48,
    G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64,
    G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80,
    G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140,
    G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184,
    G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
    G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210,
    G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245,
    G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
    G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273,
    G274, G275, G276, G277, G278, G279, G452, G483, G543, G559, G567, G651,
    G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966,
    G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078,
    G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435,
    G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3,
    G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24,
    G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44,
    G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62,
    G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78,
    G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94,
    G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138,
    G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196,
    G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208,
    G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243,
    G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255,
    G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271,
    G272, G273, G274, G275, G276, G277, G278, G279, G452, G483, G543, G559,
    G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961,
    G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072,
    G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430,
    G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n383_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n477_, new_n479_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n523_, new_n526_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT0), .B(G1083), .ZN(G367));
  XOR2_X1   g005(.A(KEYINPUT1), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  INV_X1    g010(.A(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT3), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(G223));
  NAND3_X1  g021(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n383_));
  XOR2_X1   g022(.A(new_n383_), .B(KEYINPUT4), .Z(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n386_));
  XOR2_X1   g025(.A(new_n386_), .B(KEYINPUT5), .Z(new_n387_));
  INV_X1    g026(.A(new_n387_), .ZN(new_n388_));
  NAND4_X1  g027(.A1(G44), .A2(G82), .A3(G96), .A4(G132), .ZN(new_n389_));
  XNOR2_X1  g028(.A(new_n389_), .B(KEYINPUT6), .ZN(new_n390_));
  INV_X1    g029(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g030(.A1(new_n388_), .A2(new_n391_), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n388_), .A2(G567), .B1(G2106), .B2(new_n391_), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT8), .A2(G2104), .ZN(new_n395_));
  NOR2_X1   g034(.A1(KEYINPUT8), .A2(G2104), .ZN(new_n396_));
  NOR2_X1   g035(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g036(.A1(G125), .A2(G2105), .ZN(new_n398_));
  INV_X1    g037(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g038(.A(KEYINPUT9), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g039(.A(KEYINPUT9), .ZN(new_n401_));
  NOR4_X1   g040(.A1(new_n395_), .A2(new_n396_), .A3(new_n398_), .A4(new_n401_), .ZN(new_n402_));
  NOR2_X1   g041(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g042(.A(G2105), .ZN(new_n404_));
  NAND2_X1  g043(.A1(new_n404_), .A2(KEYINPUT7), .ZN(new_n405_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n406_));
  NAND2_X1  g045(.A1(new_n406_), .A2(G2105), .ZN(new_n407_));
  NAND4_X1  g046(.A1(new_n405_), .A2(new_n407_), .A3(G101), .A4(G2104), .ZN(new_n408_));
  NAND3_X1  g047(.A1(G113), .A2(G2104), .A3(G2105), .ZN(new_n409_));
  OR2_X1    g048(.A1(KEYINPUT8), .A2(G2104), .ZN(new_n410_));
  NAND2_X1  g049(.A1(KEYINPUT8), .A2(G2104), .ZN(new_n411_));
  NAND4_X1  g050(.A1(new_n410_), .A2(new_n405_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g051(.A(G137), .ZN(new_n413_));
  OAI211_X1 g052(.A(new_n408_), .B(new_n409_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g053(.A1(new_n403_), .A2(new_n414_), .ZN(G160));
  AOI22_X1  g054(.A1(new_n397_), .A2(G124), .B1(G112), .B2(G2104), .ZN(new_n416_));
  NOR2_X1   g055(.A1(new_n416_), .A2(new_n404_), .ZN(new_n417_));
  XNOR2_X1  g056(.A(KEYINPUT7), .B(G2105), .ZN(new_n418_));
  NAND2_X1  g057(.A1(new_n418_), .A2(G2104), .ZN(new_n419_));
  INV_X1    g058(.A(G100), .ZN(new_n420_));
  INV_X1    g059(.A(G136), .ZN(new_n421_));
  OAI22_X1  g060(.A1(new_n419_), .A2(new_n420_), .B1(new_n412_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g061(.A1(new_n417_), .A2(new_n422_), .ZN(G162));
  NAND3_X1  g062(.A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n424_));
  INV_X1    g063(.A(new_n424_), .ZN(new_n425_));
  AND4_X1   g064(.A1(new_n410_), .A2(new_n405_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n426_));
  AOI21_X1  g065(.A(new_n425_), .B1(new_n426_), .B2(G138), .ZN(new_n427_));
  NAND4_X1  g066(.A1(new_n405_), .A2(new_n407_), .A3(G102), .A4(G2104), .ZN(new_n428_));
  NAND2_X1  g067(.A1(new_n428_), .A2(KEYINPUT10), .ZN(new_n429_));
  INV_X1    g068(.A(KEYINPUT10), .ZN(new_n430_));
  NAND4_X1  g069(.A1(new_n418_), .A2(new_n430_), .A3(G102), .A4(G2104), .ZN(new_n431_));
  NAND2_X1  g070(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n433_));
  NAND3_X1  g072(.A1(new_n410_), .A2(new_n411_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g073(.A(KEYINPUT11), .ZN(new_n435_));
  NAND2_X1  g074(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g075(.A1(new_n397_), .A2(KEYINPUT11), .A3(new_n433_), .ZN(new_n437_));
  NAND2_X1  g076(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g077(.A1(new_n427_), .A2(new_n432_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g078(.A(new_n439_), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n441_));
  INV_X1    g080(.A(G543), .ZN(new_n442_));
  AOI21_X1  g081(.A(new_n441_), .B1(G62), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g082(.A(G75), .ZN(new_n444_));
  OAI21_X1  g083(.A(new_n443_), .B1(new_n444_), .B2(new_n442_), .ZN(new_n445_));
  AOI21_X1  g084(.A(G651), .B1(new_n442_), .B2(G88), .ZN(new_n446_));
  INV_X1    g085(.A(G50), .ZN(new_n447_));
  OAI21_X1  g086(.A(new_n446_), .B1(new_n447_), .B2(new_n442_), .ZN(new_n448_));
  NAND2_X1  g087(.A1(new_n445_), .A2(new_n448_), .ZN(G166));
  NAND2_X1  g088(.A1(G76), .A2(G543), .ZN(new_n450_));
  INV_X1    g089(.A(G63), .ZN(new_n451_));
  OAI211_X1 g090(.A(new_n450_), .B(G651), .C1(new_n451_), .C2(G543), .ZN(new_n452_));
  NAND2_X1  g091(.A1(G51), .A2(G543), .ZN(new_n453_));
  INV_X1    g092(.A(G89), .ZN(new_n454_));
  OAI211_X1 g093(.A(new_n453_), .B(new_n441_), .C1(new_n454_), .C2(G543), .ZN(new_n455_));
  NAND2_X1  g094(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n457_));
  XNOR2_X1  g096(.A(new_n456_), .B(new_n457_), .ZN(G168));
  NAND3_X1  g097(.A1(G77), .A2(G543), .A3(G651), .ZN(new_n459_));
  XOR2_X1   g098(.A(new_n459_), .B(KEYINPUT14), .Z(new_n460_));
  NAND3_X1  g099(.A1(new_n442_), .A2(G64), .A3(G651), .ZN(new_n461_));
  XNOR2_X1  g100(.A(new_n461_), .B(KEYINPUT13), .ZN(new_n462_));
  OR2_X1    g101(.A1(G90), .A2(G543), .ZN(new_n463_));
  OAI211_X1 g102(.A(new_n463_), .B(new_n441_), .C1(G52), .C2(new_n442_), .ZN(new_n464_));
  NAND3_X1  g103(.A1(new_n460_), .A2(new_n462_), .A3(new_n464_), .ZN(G301));
  XOR2_X1   g104(.A(G301), .B(KEYINPUT15), .Z(G171));
  NAND3_X1  g105(.A1(new_n441_), .A2(G43), .A3(G543), .ZN(new_n467_));
  INV_X1    g106(.A(KEYINPUT16), .ZN(new_n468_));
  XNOR2_X1  g107(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  OR2_X1    g108(.A1(G56), .A2(G543), .ZN(new_n470_));
  OAI211_X1 g109(.A(new_n470_), .B(G651), .C1(G68), .C2(new_n442_), .ZN(new_n471_));
  NOR2_X1   g110(.A1(G543), .A2(G651), .ZN(new_n472_));
  NAND2_X1  g111(.A1(new_n472_), .A2(G81), .ZN(new_n473_));
  NAND3_X1  g112(.A1(new_n469_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g113(.A(G860), .ZN(new_n475_));
  OR2_X1    g114(.A1(new_n474_), .A2(new_n475_), .ZN(G153));
  AND2_X1   g115(.A1(G483), .A2(G661), .ZN(new_n477_));
  NAND3_X1  g116(.A1(G319), .A2(G36), .A3(new_n477_), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n479_));
  NAND3_X1  g118(.A1(G319), .A2(new_n477_), .A3(new_n479_), .ZN(G188));
  AOI21_X1  g119(.A(new_n441_), .B1(G65), .B2(new_n442_), .ZN(new_n481_));
  INV_X1    g120(.A(G78), .ZN(new_n482_));
  OAI21_X1  g121(.A(new_n481_), .B1(new_n482_), .B2(new_n442_), .ZN(new_n483_));
  AOI21_X1  g122(.A(G651), .B1(new_n442_), .B2(G91), .ZN(new_n484_));
  INV_X1    g123(.A(G53), .ZN(new_n485_));
  OAI21_X1  g124(.A(new_n484_), .B1(new_n485_), .B2(new_n442_), .ZN(new_n486_));
  NAND2_X1  g125(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g126(.A(new_n487_), .ZN(G299));
  XNOR2_X1  g127(.A(new_n456_), .B(KEYINPUT12), .ZN(G286));
  INV_X1    g128(.A(G166), .ZN(G303));
  AOI21_X1  g129(.A(G651), .B1(new_n442_), .B2(G87), .ZN(new_n491_));
  INV_X1    g130(.A(G49), .ZN(new_n492_));
  OAI21_X1  g131(.A(new_n491_), .B1(new_n492_), .B2(new_n442_), .ZN(new_n493_));
  OR3_X1    g132(.A1(new_n442_), .A2(new_n441_), .A3(G74), .ZN(new_n494_));
  NAND2_X1  g133(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g134(.A(new_n495_), .ZN(G288));
  INV_X1    g135(.A(G61), .ZN(new_n497_));
  OAI21_X1  g136(.A(G651), .B1(new_n497_), .B2(G543), .ZN(new_n498_));
  INV_X1    g137(.A(new_n472_), .ZN(new_n499_));
  OAI221_X1 g138(.A(new_n498_), .B1(G48), .B2(new_n442_), .C1(new_n499_), .C2(G86), .ZN(new_n500_));
  NAND3_X1  g139(.A1(G73), .A2(G543), .A3(G651), .ZN(new_n501_));
  XNOR2_X1  g140(.A(new_n501_), .B(KEYINPUT17), .ZN(new_n502_));
  NAND2_X1  g141(.A1(new_n500_), .A2(new_n502_), .ZN(G305));
  AOI21_X1  g142(.A(new_n441_), .B1(G60), .B2(new_n442_), .ZN(new_n504_));
  NAND2_X1  g143(.A1(G72), .A2(G543), .ZN(new_n505_));
  AOI21_X1  g144(.A(G651), .B1(new_n442_), .B2(G85), .ZN(new_n506_));
  NAND2_X1  g145(.A1(G47), .A2(G543), .ZN(new_n507_));
  AOI22_X1  g146(.A1(new_n504_), .A2(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(G290));
  NAND2_X1  g147(.A1(G301), .A2(G868), .ZN(new_n509_));
  AND3_X1   g148(.A1(new_n441_), .A2(G54), .A3(G543), .ZN(new_n510_));
  NAND2_X1  g149(.A1(new_n472_), .A2(G92), .ZN(new_n511_));
  INV_X1    g150(.A(G79), .ZN(new_n512_));
  NAND2_X1  g151(.A1(new_n512_), .A2(G543), .ZN(new_n513_));
  INV_X1    g152(.A(new_n513_), .ZN(new_n514_));
  OAI21_X1  g153(.A(G651), .B1(G66), .B2(G543), .ZN(new_n515_));
  OAI21_X1  g154(.A(new_n511_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g155(.A1(new_n516_), .A2(KEYINPUT18), .ZN(new_n517_));
  INV_X1    g156(.A(KEYINPUT18), .ZN(new_n518_));
  OAI211_X1 g157(.A(new_n511_), .B(new_n518_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n519_));
  AOI21_X1  g158(.A(new_n510_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g159(.A(new_n509_), .B1(new_n520_), .B2(G868), .ZN(G284));
  OAI21_X1  g160(.A(new_n509_), .B1(new_n520_), .B2(G868), .ZN(G321));
  NOR2_X1   g161(.A1(G299), .A2(G868), .ZN(new_n523_));
  AOI21_X1  g162(.A(new_n523_), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g163(.A(new_n523_), .B1(G168), .B2(G868), .ZN(G280));
  NAND2_X1  g164(.A1(new_n475_), .A2(G559), .ZN(new_n526_));
  NAND2_X1  g165(.A1(new_n520_), .A2(new_n526_), .ZN(G148));
  INV_X1    g166(.A(G868), .ZN(new_n528_));
  NAND2_X1  g167(.A1(new_n474_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g168(.A(new_n520_), .ZN(new_n530_));
  NOR2_X1   g169(.A1(new_n530_), .A2(G559), .ZN(new_n531_));
  OAI21_X1  g170(.A(new_n529_), .B1(new_n531_), .B2(new_n528_), .ZN(G282));
  OAI21_X1  g171(.A(new_n529_), .B1(new_n531_), .B2(new_n528_), .ZN(G323));
  NAND2_X1  g172(.A1(G111), .A2(G2104), .ZN(new_n534_));
  NAND2_X1  g173(.A1(new_n410_), .A2(new_n411_), .ZN(new_n535_));
  INV_X1    g174(.A(G123), .ZN(new_n536_));
  OAI21_X1  g175(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  AND2_X1   g176(.A1(new_n418_), .A2(G2104), .ZN(new_n538_));
  AOI22_X1  g177(.A1(G2105), .A2(new_n537_), .B1(new_n538_), .B2(G99), .ZN(new_n539_));
  NAND3_X1  g178(.A1(new_n426_), .A2(KEYINPUT19), .A3(G135), .ZN(new_n540_));
  INV_X1    g179(.A(KEYINPUT19), .ZN(new_n541_));
  INV_X1    g180(.A(G135), .ZN(new_n542_));
  OAI21_X1  g181(.A(new_n541_), .B1(new_n412_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g182(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g183(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  OR2_X1    g184(.A1(new_n545_), .A2(G2096), .ZN(new_n546_));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n547_));
  OAI21_X1  g186(.A(new_n547_), .B1(new_n397_), .B2(G2105), .ZN(new_n548_));
  NAND3_X1  g187(.A1(new_n535_), .A2(KEYINPUT20), .A3(new_n404_), .ZN(new_n549_));
  NAND3_X1  g188(.A1(new_n548_), .A2(new_n538_), .A3(new_n549_), .ZN(new_n550_));
  XOR2_X1   g189(.A(new_n550_), .B(G2100), .Z(new_n551_));
  NAND2_X1  g190(.A1(new_n545_), .A2(G2096), .ZN(new_n552_));
  NAND3_X1  g191(.A1(new_n546_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  XOR2_X1   g192(.A(new_n553_), .B(KEYINPUT21), .Z(G156));
  XOR2_X1   g193(.A(G2451), .B(G2454), .Z(new_n555_));
  XNOR2_X1  g194(.A(new_n555_), .B(KEYINPUT24), .ZN(new_n556_));
  XOR2_X1   g195(.A(G2443), .B(G2446), .Z(new_n557_));
  XNOR2_X1  g196(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g197(.A(KEYINPUT22), .ZN(new_n559_));
  XNOR2_X1  g198(.A(KEYINPUT23), .B(G2435), .ZN(new_n560_));
  XNOR2_X1  g199(.A(new_n560_), .B(G2438), .ZN(new_n561_));
  XNOR2_X1  g200(.A(G2427), .B(G2430), .ZN(new_n562_));
  AOI21_X1  g201(.A(new_n559_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g202(.A(new_n563_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n564_));
  XNOR2_X1  g203(.A(new_n558_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n566_));
  INV_X1    g205(.A(new_n566_), .ZN(new_n567_));
  OR2_X1    g206(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g207(.A1(new_n565_), .A2(new_n567_), .ZN(new_n569_));
  AND3_X1   g208(.A1(new_n568_), .A2(G14), .A3(new_n569_), .ZN(G401));
  XNOR2_X1  g209(.A(G2084), .B(G2090), .ZN(new_n571_));
  XNOR2_X1  g210(.A(G2096), .B(G2100), .ZN(new_n572_));
  XNOR2_X1  g211(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g212(.A(G2072), .B(G2078), .ZN(new_n574_));
  XNOR2_X1  g213(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n576_));
  XNOR2_X1  g215(.A(new_n576_), .B(KEYINPUT25), .ZN(new_n577_));
  XNOR2_X1  g216(.A(new_n577_), .B(KEYINPUT26), .ZN(new_n578_));
  XNOR2_X1  g217(.A(new_n575_), .B(new_n578_), .ZN(G227));
  XOR2_X1   g218(.A(G1971), .B(G1976), .Z(new_n580_));
  INV_X1    g219(.A(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g220(.A(G1956), .B(G2474), .ZN(new_n582_));
  XNOR2_X1  g221(.A(G1961), .B(G1966), .ZN(new_n583_));
  NOR3_X1   g222(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g223(.A(new_n584_), .B(KEYINPUT27), .ZN(new_n585_));
  NAND3_X1  g224(.A1(new_n580_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n586_));
  AND2_X1   g225(.A1(new_n582_), .A2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g226(.A(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n588_));
  OAI211_X1 g227(.A(new_n585_), .B(new_n586_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g228(.A(new_n589_), .B(G1991), .ZN(new_n590_));
  XNOR2_X1  g229(.A(G1981), .B(G1986), .ZN(new_n591_));
  XNOR2_X1  g230(.A(new_n591_), .B(KEYINPUT28), .ZN(new_n592_));
  XNOR2_X1  g231(.A(new_n592_), .B(G1996), .ZN(new_n593_));
  INV_X1    g232(.A(new_n593_), .ZN(new_n594_));
  OR2_X1    g233(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g234(.A1(new_n590_), .A2(new_n594_), .ZN(new_n596_));
  NAND2_X1  g235(.A1(new_n595_), .A2(new_n596_), .ZN(G229));
  NAND2_X1  g236(.A1(G162), .A2(G29), .ZN(new_n598_));
  OAI21_X1  g237(.A(new_n598_), .B1(G29), .B2(G35), .ZN(new_n599_));
  INV_X1    g238(.A(G2090), .ZN(new_n600_));
  OR2_X1    g239(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g240(.A1(G16), .A2(G22), .ZN(new_n602_));
  AOI21_X1  g241(.A(new_n602_), .B1(G166), .B2(G16), .ZN(new_n603_));
  AND2_X1   g242(.A1(new_n603_), .A2(G1971), .ZN(new_n604_));
  NOR2_X1   g243(.A1(new_n603_), .A2(G1971), .ZN(new_n605_));
  AND3_X1   g244(.A1(KEYINPUT35), .A2(G11), .A3(G868), .ZN(new_n606_));
  OAI22_X1  g245(.A1(KEYINPUT35), .A2(G11), .B1(G28), .B2(G29), .ZN(new_n607_));
  NOR4_X1   g246(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  INV_X1    g247(.A(G301), .ZN(new_n609_));
  NAND2_X1  g248(.A1(new_n609_), .A2(G16), .ZN(new_n610_));
  OAI21_X1  g249(.A(new_n610_), .B1(G5), .B2(G16), .ZN(new_n611_));
  INV_X1    g250(.A(G1961), .ZN(new_n612_));
  NAND2_X1  g251(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g252(.A1(G16), .A2(G21), .ZN(new_n614_));
  AOI21_X1  g253(.A(new_n614_), .B1(G168), .B2(G16), .ZN(new_n615_));
  NAND2_X1  g254(.A1(new_n615_), .A2(G1966), .ZN(new_n616_));
  NAND4_X1  g255(.A1(new_n601_), .A2(new_n608_), .A3(new_n613_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g256(.A1(new_n599_), .A2(new_n600_), .ZN(new_n618_));
  OAI221_X1 g257(.A(new_n618_), .B1(new_n612_), .B2(new_n611_), .C1(G1966), .C2(new_n615_), .ZN(new_n619_));
  NOR2_X1   g258(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g259(.A(G16), .ZN(new_n621_));
  INV_X1    g260(.A(G23), .ZN(new_n622_));
  AND2_X1   g261(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n623_));
  NOR2_X1   g262(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n624_));
  OAI21_X1  g263(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n626_));
  OR2_X1    g265(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g266(.A1(new_n625_), .A2(new_n626_), .ZN(new_n628_));
  OAI211_X1 g267(.A(new_n627_), .B(new_n628_), .C1(new_n621_), .C2(new_n495_), .ZN(new_n629_));
  INV_X1    g268(.A(G1976), .ZN(new_n630_));
  XNOR2_X1  g269(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n632_));
  OR2_X1    g271(.A1(new_n632_), .A2(G1981), .ZN(new_n633_));
  NOR2_X1   g272(.A1(G16), .A2(G20), .ZN(new_n634_));
  AOI21_X1  g273(.A(new_n634_), .B1(new_n487_), .B2(G16), .ZN(new_n635_));
  XOR2_X1   g274(.A(new_n635_), .B(G1956), .Z(new_n636_));
  NAND2_X1  g275(.A1(new_n632_), .A2(G1981), .ZN(new_n637_));
  NAND4_X1  g276(.A1(new_n631_), .A2(new_n633_), .A3(new_n636_), .A4(new_n637_), .ZN(new_n638_));
  MUX2_X1   g277(.A(G19), .B(new_n474_), .S(G16), .Z(new_n639_));
  NAND2_X1  g278(.A1(new_n639_), .A2(G1341), .ZN(new_n640_));
  INV_X1    g279(.A(G29), .ZN(new_n641_));
  OAI21_X1  g280(.A(new_n640_), .B1(new_n641_), .B2(new_n545_), .ZN(new_n642_));
  MUX2_X1   g281(.A(G24), .B(G290), .S(G16), .Z(new_n643_));
  XNOR2_X1  g282(.A(new_n643_), .B(G1986), .ZN(new_n644_));
  NOR2_X1   g283(.A1(new_n639_), .A2(G1341), .ZN(new_n645_));
  NOR4_X1   g284(.A1(new_n638_), .A2(new_n642_), .A3(new_n644_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g285(.A(G103), .ZN(new_n647_));
  INV_X1    g286(.A(G139), .ZN(new_n648_));
  OAI22_X1  g287(.A1(new_n419_), .A2(new_n647_), .B1(new_n412_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g288(.A1(new_n397_), .A2(G127), .ZN(new_n650_));
  NAND2_X1  g289(.A1(G115), .A2(G2104), .ZN(new_n651_));
  AOI21_X1  g290(.A(new_n404_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g291(.A(G29), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g292(.A1(new_n641_), .A2(G33), .ZN(new_n654_));
  XNOR2_X1  g293(.A(new_n654_), .B(KEYINPUT30), .ZN(new_n655_));
  NAND2_X1  g294(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g295(.A(new_n656_), .B(G2072), .ZN(new_n657_));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n658_));
  AOI21_X1  g297(.A(new_n658_), .B1(new_n520_), .B2(G16), .ZN(new_n659_));
  AOI21_X1  g298(.A(new_n657_), .B1(G1348), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g299(.A1(new_n620_), .A2(new_n646_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g300(.A1(new_n641_), .A2(G27), .ZN(new_n662_));
  OAI21_X1  g301(.A(new_n662_), .B1(G164), .B2(new_n641_), .ZN(new_n663_));
  XNOR2_X1  g302(.A(new_n663_), .B(G2078), .ZN(new_n664_));
  OR2_X1    g303(.A1(new_n664_), .A2(KEYINPUT34), .ZN(new_n665_));
  NOR2_X1   g304(.A1(G25), .A2(G29), .ZN(new_n666_));
  AOI22_X1  g305(.A1(new_n397_), .A2(G119), .B1(G107), .B2(G2104), .ZN(new_n667_));
  NOR2_X1   g306(.A1(new_n667_), .A2(new_n404_), .ZN(new_n668_));
  INV_X1    g307(.A(G95), .ZN(new_n669_));
  INV_X1    g308(.A(G131), .ZN(new_n670_));
  OAI22_X1  g309(.A1(new_n419_), .A2(new_n669_), .B1(new_n412_), .B2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g310(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g311(.A(new_n666_), .B1(new_n672_), .B2(G29), .ZN(new_n673_));
  XNOR2_X1  g312(.A(KEYINPUT38), .B(G1991), .ZN(new_n674_));
  XOR2_X1   g313(.A(new_n673_), .B(new_n674_), .Z(new_n675_));
  NAND2_X1  g314(.A1(new_n641_), .A2(G32), .ZN(new_n676_));
  NAND2_X1  g315(.A1(new_n397_), .A2(G2105), .ZN(new_n677_));
  INV_X1    g316(.A(G129), .ZN(new_n678_));
  INV_X1    g317(.A(G141), .ZN(new_n679_));
  OAI22_X1  g318(.A1(new_n677_), .A2(new_n678_), .B1(new_n412_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n681_));
  XNOR2_X1  g320(.A(new_n681_), .B(KEYINPUT31), .ZN(new_n682_));
  INV_X1    g321(.A(G105), .ZN(new_n683_));
  OAI21_X1  g322(.A(new_n682_), .B1(new_n419_), .B2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g323(.A1(new_n680_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g324(.A(new_n676_), .B1(new_n685_), .B2(new_n641_), .ZN(new_n686_));
  XNOR2_X1  g325(.A(new_n686_), .B(G1996), .ZN(new_n687_));
  NOR2_X1   g326(.A1(new_n659_), .A2(G1348), .ZN(new_n688_));
  NOR3_X1   g327(.A1(new_n675_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g328(.A1(new_n664_), .A2(KEYINPUT34), .ZN(new_n690_));
  NAND3_X1  g329(.A1(new_n665_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  AOI22_X1  g330(.A1(new_n538_), .A2(G104), .B1(new_n426_), .B2(G140), .ZN(new_n692_));
  NOR2_X1   g331(.A1(new_n535_), .A2(new_n404_), .ZN(new_n693_));
  NAND2_X1  g332(.A1(new_n693_), .A2(G128), .ZN(new_n694_));
  NAND3_X1  g333(.A1(G116), .A2(G2104), .A3(G2105), .ZN(new_n695_));
  INV_X1    g334(.A(KEYINPUT32), .ZN(new_n696_));
  XNOR2_X1  g335(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  NAND4_X1  g336(.A1(new_n692_), .A2(KEYINPUT33), .A3(new_n694_), .A4(new_n697_), .ZN(new_n698_));
  INV_X1    g337(.A(KEYINPUT33), .ZN(new_n699_));
  INV_X1    g338(.A(G104), .ZN(new_n700_));
  INV_X1    g339(.A(G140), .ZN(new_n701_));
  OAI22_X1  g340(.A1(new_n419_), .A2(new_n700_), .B1(new_n412_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g341(.A(G128), .ZN(new_n703_));
  OAI21_X1  g342(.A(new_n697_), .B1(new_n677_), .B2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g343(.A(new_n699_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  AND2_X1   g344(.A1(new_n698_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g345(.A1(new_n706_), .A2(G29), .ZN(new_n707_));
  OAI21_X1  g346(.A(new_n707_), .B1(G26), .B2(G29), .ZN(new_n708_));
  INV_X1    g347(.A(G2067), .ZN(new_n709_));
  OR2_X1    g348(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g349(.A1(new_n708_), .A2(new_n709_), .ZN(new_n711_));
  INV_X1    g350(.A(G34), .ZN(new_n712_));
  AND2_X1   g351(.A1(new_n712_), .A2(KEYINPUT29), .ZN(new_n713_));
  NOR2_X1   g352(.A1(new_n712_), .A2(KEYINPUT29), .ZN(new_n714_));
  OAI21_X1  g353(.A(new_n641_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g354(.A(new_n715_), .B1(G160), .B2(new_n641_), .ZN(new_n716_));
  XOR2_X1   g355(.A(new_n716_), .B(G2084), .Z(new_n717_));
  NAND3_X1  g356(.A1(new_n710_), .A2(new_n711_), .A3(new_n717_), .ZN(new_n718_));
  NOR3_X1   g357(.A1(new_n661_), .A2(new_n691_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g358(.A(KEYINPUT39), .ZN(new_n720_));
  XNOR2_X1  g359(.A(new_n719_), .B(new_n720_), .ZN(G311));
  XNOR2_X1  g360(.A(new_n719_), .B(KEYINPUT39), .ZN(G150));
  OAI21_X1  g361(.A(G153), .B1(new_n530_), .B2(new_n526_), .ZN(new_n723_));
  NAND3_X1  g362(.A1(new_n441_), .A2(G55), .A3(G543), .ZN(new_n724_));
  XNOR2_X1  g363(.A(new_n724_), .B(KEYINPUT40), .ZN(new_n725_));
  OR2_X1    g364(.A1(new_n442_), .A2(G80), .ZN(new_n726_));
  OAI21_X1  g365(.A(G651), .B1(G67), .B2(G543), .ZN(new_n727_));
  INV_X1    g366(.A(new_n727_), .ZN(new_n728_));
  AOI22_X1  g367(.A1(new_n726_), .A2(new_n728_), .B1(G93), .B2(new_n472_), .ZN(new_n729_));
  NAND2_X1  g368(.A1(new_n725_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g369(.A(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g370(.A(new_n731_), .B(new_n474_), .ZN(new_n732_));
  XNOR2_X1  g371(.A(new_n723_), .B(new_n732_), .ZN(G145));
  XOR2_X1   g372(.A(KEYINPUT44), .B(G37), .Z(new_n734_));
  INV_X1    g373(.A(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g374(.A(new_n550_), .B(KEYINPUT43), .ZN(new_n736_));
  NAND2_X1  g375(.A1(new_n736_), .A2(new_n545_), .ZN(new_n737_));
  INV_X1    g376(.A(KEYINPUT43), .ZN(new_n738_));
  XNOR2_X1  g377(.A(new_n550_), .B(new_n738_), .ZN(new_n739_));
  INV_X1    g378(.A(new_n545_), .ZN(new_n740_));
  NAND2_X1  g379(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g380(.A1(new_n737_), .A2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g381(.A(G162), .B1(new_n403_), .B2(new_n414_), .ZN(new_n743_));
  OAI21_X1  g382(.A(G160), .B1(new_n417_), .B2(new_n422_), .ZN(new_n744_));
  NAND2_X1  g383(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g384(.A(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g385(.A(new_n742_), .B(new_n746_), .ZN(new_n747_));
  NAND2_X1  g386(.A1(new_n698_), .A2(new_n705_), .ZN(new_n748_));
  NAND2_X1  g387(.A1(new_n748_), .A2(new_n685_), .ZN(new_n749_));
  OR2_X1    g388(.A1(new_n680_), .A2(new_n684_), .ZN(new_n750_));
  NAND3_X1  g389(.A1(new_n698_), .A2(new_n750_), .A3(new_n705_), .ZN(new_n751_));
  OAI21_X1  g390(.A(KEYINPUT41), .B1(new_n649_), .B2(new_n652_), .ZN(new_n752_));
  NAND2_X1  g391(.A1(new_n650_), .A2(new_n651_), .ZN(new_n753_));
  NAND2_X1  g392(.A1(new_n753_), .A2(G2105), .ZN(new_n754_));
  INV_X1    g393(.A(KEYINPUT41), .ZN(new_n755_));
  NAND2_X1  g394(.A1(new_n426_), .A2(G139), .ZN(new_n756_));
  NAND2_X1  g395(.A1(new_n538_), .A2(G103), .ZN(new_n757_));
  NAND4_X1  g396(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .A4(new_n757_), .ZN(new_n758_));
  NAND3_X1  g397(.A1(G164), .A2(new_n752_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g398(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g399(.A(G164), .B1(new_n752_), .B2(new_n758_), .ZN(new_n761_));
  OAI211_X1 g400(.A(new_n749_), .B(new_n751_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g401(.A1(new_n758_), .A2(new_n752_), .ZN(new_n763_));
  NAND2_X1  g402(.A1(new_n763_), .A2(new_n439_), .ZN(new_n764_));
  AND3_X1   g403(.A1(new_n698_), .A2(new_n750_), .A3(new_n705_), .ZN(new_n765_));
  AOI21_X1  g404(.A(new_n750_), .B1(new_n698_), .B2(new_n705_), .ZN(new_n766_));
  OAI211_X1 g405(.A(new_n759_), .B(new_n764_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g406(.A1(new_n693_), .A2(G130), .ZN(new_n768_));
  XOR2_X1   g407(.A(new_n768_), .B(KEYINPUT42), .Z(new_n769_));
  INV_X1    g408(.A(new_n672_), .ZN(new_n770_));
  NAND2_X1  g409(.A1(new_n538_), .A2(G106), .ZN(new_n771_));
  NAND2_X1  g410(.A1(new_n426_), .A2(G142), .ZN(new_n772_));
  NAND3_X1  g411(.A1(G118), .A2(G2104), .A3(G2105), .ZN(new_n773_));
  NAND3_X1  g412(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g413(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g414(.A1(new_n769_), .A2(new_n770_), .A3(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g415(.A(new_n768_), .B(KEYINPUT42), .ZN(new_n777_));
  OAI21_X1  g416(.A(new_n672_), .B1(new_n777_), .B2(new_n774_), .ZN(new_n778_));
  AND2_X1   g417(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  AND3_X1   g418(.A1(new_n762_), .A2(new_n767_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g419(.A(new_n779_), .B1(new_n762_), .B2(new_n767_), .ZN(new_n781_));
  OAI21_X1  g420(.A(new_n747_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g421(.A1(new_n762_), .A2(new_n767_), .ZN(new_n783_));
  INV_X1    g422(.A(new_n779_), .ZN(new_n784_));
  NAND2_X1  g423(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g424(.A(new_n742_), .B(new_n745_), .ZN(new_n786_));
  NAND3_X1  g425(.A1(new_n762_), .A2(new_n767_), .A3(new_n779_), .ZN(new_n787_));
  NAND3_X1  g426(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g427(.A(new_n735_), .B1(new_n782_), .B2(new_n788_), .ZN(G395));
  INV_X1    g428(.A(KEYINPUT45), .ZN(new_n790_));
  XNOR2_X1  g429(.A(new_n520_), .B(new_n487_), .ZN(new_n791_));
  OR2_X1    g430(.A1(new_n791_), .A2(new_n732_), .ZN(new_n792_));
  NAND2_X1  g431(.A1(new_n791_), .A2(new_n732_), .ZN(new_n793_));
  AOI21_X1  g432(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g433(.A(new_n531_), .ZN(new_n795_));
  NAND2_X1  g434(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g435(.A(new_n795_), .B1(new_n792_), .B2(new_n790_), .ZN(new_n797_));
  INV_X1    g436(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g437(.A(new_n796_), .B1(new_n798_), .B2(new_n794_), .ZN(new_n799_));
  XNOR2_X1  g438(.A(G305), .B(G288), .ZN(new_n800_));
  XNOR2_X1  g439(.A(G166), .B(G290), .ZN(new_n801_));
  XOR2_X1   g440(.A(new_n800_), .B(new_n801_), .Z(new_n802_));
  INV_X1    g441(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g442(.A1(new_n799_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g443(.A(new_n796_), .B(new_n802_), .C1(new_n798_), .C2(new_n794_), .ZN(new_n805_));
  AOI21_X1  g444(.A(new_n528_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g445(.A1(new_n731_), .A2(G868), .ZN(new_n807_));
  OAI21_X1  g446(.A(KEYINPUT46), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g447(.A(new_n805_), .ZN(new_n809_));
  AND2_X1   g448(.A1(new_n792_), .A2(new_n793_), .ZN(new_n810_));
  OAI21_X1  g449(.A(new_n797_), .B1(new_n810_), .B2(new_n790_), .ZN(new_n811_));
  AOI21_X1  g450(.A(new_n802_), .B1(new_n811_), .B2(new_n796_), .ZN(new_n812_));
  OAI21_X1  g451(.A(G868), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g452(.A(KEYINPUT46), .ZN(new_n814_));
  INV_X1    g453(.A(new_n807_), .ZN(new_n815_));
  NAND3_X1  g454(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g455(.A1(new_n808_), .A2(new_n816_), .ZN(G295));
  NAND2_X1  g456(.A1(new_n813_), .A2(new_n815_), .ZN(G331));
  XNOR2_X1  g457(.A(G286), .B(G301), .ZN(new_n819_));
  NAND2_X1  g458(.A1(new_n810_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g459(.A1(new_n792_), .A2(new_n793_), .ZN(new_n821_));
  INV_X1    g460(.A(new_n819_), .ZN(new_n822_));
  NAND2_X1  g461(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND3_X1   g462(.A1(new_n820_), .A2(new_n803_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g463(.A(new_n803_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n825_));
  OAI21_X1  g464(.A(new_n734_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g465(.A(new_n826_), .ZN(G397));
  INV_X1    g466(.A(G1384), .ZN(new_n828_));
  NAND3_X1  g467(.A1(new_n397_), .A2(new_n418_), .A3(G138), .ZN(new_n829_));
  AOI21_X1  g468(.A(KEYINPUT11), .B1(new_n397_), .B2(new_n433_), .ZN(new_n830_));
  AND4_X1   g469(.A1(KEYINPUT11), .A2(new_n410_), .A3(new_n411_), .A4(new_n433_), .ZN(new_n831_));
  OAI211_X1 g470(.A(new_n829_), .B(new_n424_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n832_));
  AND2_X1   g471(.A1(new_n429_), .A2(new_n431_), .ZN(new_n833_));
  OAI21_X1  g472(.A(new_n828_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g473(.A(new_n834_), .ZN(new_n835_));
  NAND3_X1  g474(.A1(new_n410_), .A2(new_n399_), .A3(new_n411_), .ZN(new_n836_));
  XNOR2_X1  g475(.A(new_n836_), .B(new_n401_), .ZN(new_n837_));
  INV_X1    g476(.A(new_n409_), .ZN(new_n838_));
  AOI21_X1  g477(.A(new_n838_), .B1(new_n426_), .B2(G137), .ZN(new_n839_));
  NAND4_X1  g478(.A1(new_n837_), .A2(new_n839_), .A3(G40), .A4(new_n408_), .ZN(new_n840_));
  NOR2_X1   g479(.A1(new_n835_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g480(.A1(new_n841_), .A2(new_n706_), .A3(new_n709_), .ZN(new_n842_));
  NOR2_X1   g481(.A1(new_n842_), .A2(KEYINPUT50), .ZN(new_n843_));
  INV_X1    g482(.A(KEYINPUT50), .ZN(new_n844_));
  NOR2_X1   g483(.A1(new_n750_), .A2(G1996), .ZN(new_n845_));
  NAND2_X1  g484(.A1(new_n841_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g485(.A1(new_n706_), .A2(new_n709_), .ZN(new_n847_));
  OAI21_X1  g486(.A(new_n844_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g487(.A(new_n843_), .B1(new_n848_), .B2(new_n842_), .ZN(new_n849_));
  NAND2_X1  g488(.A1(new_n841_), .A2(G290), .ZN(new_n850_));
  XOR2_X1   g489(.A(new_n850_), .B(KEYINPUT48), .Z(new_n851_));
  XOR2_X1   g490(.A(KEYINPUT47), .B(G1986), .Z(new_n852_));
  NAND2_X1  g491(.A1(new_n841_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g492(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g493(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g494(.A1(new_n847_), .A2(new_n841_), .ZN(new_n856_));
  AND2_X1   g495(.A1(new_n750_), .A2(G1996), .ZN(new_n857_));
  OAI21_X1  g496(.A(new_n841_), .B1(new_n857_), .B2(new_n845_), .ZN(new_n858_));
  AND3_X1   g497(.A1(new_n856_), .A2(new_n858_), .A3(new_n842_), .ZN(new_n859_));
  AND2_X1   g498(.A1(new_n672_), .A2(new_n674_), .ZN(new_n860_));
  NOR2_X1   g499(.A1(new_n672_), .A2(new_n674_), .ZN(new_n861_));
  OAI21_X1  g500(.A(new_n841_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g501(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g502(.A(new_n849_), .B1(new_n855_), .B2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g503(.A1(new_n859_), .A2(new_n841_), .A3(new_n860_), .ZN(new_n865_));
  NAND2_X1  g504(.A1(new_n865_), .A2(KEYINPUT49), .ZN(new_n866_));
  OR2_X1    g505(.A1(new_n865_), .A2(KEYINPUT49), .ZN(new_n867_));
  AOI21_X1  g506(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g507(.A(G8), .ZN(new_n869_));
  INV_X1    g508(.A(G1981), .ZN(new_n870_));
  NAND3_X1  g509(.A1(new_n500_), .A2(new_n502_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g510(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g511(.A(new_n870_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n873_));
  OAI21_X1  g512(.A(KEYINPUT51), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g513(.A1(G305), .A2(G1981), .ZN(new_n875_));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n876_));
  NAND3_X1  g515(.A1(new_n875_), .A2(new_n876_), .A3(new_n871_), .ZN(new_n877_));
  NAND2_X1  g516(.A1(new_n874_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g517(.A1(G288), .A2(G1976), .ZN(new_n879_));
  AOI21_X1  g518(.A(new_n872_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g519(.A(G40), .ZN(new_n881_));
  NOR3_X1   g520(.A1(new_n403_), .A2(new_n414_), .A3(new_n881_), .ZN(new_n882_));
  AOI211_X1 g521(.A(new_n869_), .B(new_n880_), .C1(new_n835_), .C2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g522(.A1(new_n495_), .A2(G1976), .ZN(new_n884_));
  OAI211_X1 g523(.A(G8), .B(new_n884_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n885_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n886_));
  NAND2_X1  g525(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g526(.A1(new_n882_), .A2(new_n828_), .A3(new_n439_), .ZN(new_n888_));
  NAND4_X1  g527(.A1(new_n888_), .A2(G8), .A3(new_n874_), .A4(new_n877_), .ZN(new_n889_));
  AOI21_X1  g528(.A(new_n886_), .B1(G288), .B2(new_n630_), .ZN(new_n890_));
  NAND4_X1  g529(.A1(new_n888_), .A2(G8), .A3(new_n884_), .A4(new_n890_), .ZN(new_n891_));
  NAND3_X1  g530(.A1(new_n887_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  OAI21_X1  g531(.A(G1971), .B1(new_n834_), .B2(new_n840_), .ZN(new_n893_));
  NAND4_X1  g532(.A1(new_n882_), .A2(new_n828_), .A3(G2090), .A4(new_n439_), .ZN(new_n894_));
  AOI211_X1 g533(.A(new_n869_), .B(G166), .C1(new_n893_), .C2(new_n894_), .ZN(new_n895_));
  AND4_X1   g534(.A1(G8), .A2(new_n893_), .A3(G166), .A4(new_n894_), .ZN(new_n896_));
  NOR3_X1   g535(.A1(new_n892_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  OAI21_X1  g536(.A(G1966), .B1(new_n834_), .B2(new_n840_), .ZN(new_n898_));
  OAI21_X1  g537(.A(KEYINPUT52), .B1(G168), .B2(new_n869_), .ZN(new_n899_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n900_));
  NAND3_X1  g539(.A1(G286), .A2(new_n900_), .A3(G8), .ZN(new_n901_));
  NAND2_X1  g540(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  NAND4_X1  g541(.A1(new_n882_), .A2(new_n828_), .A3(G2084), .A4(new_n439_), .ZN(new_n903_));
  AND4_X1   g542(.A1(G8), .A2(new_n898_), .A3(new_n902_), .A4(new_n903_), .ZN(new_n904_));
  AOI21_X1  g543(.A(new_n883_), .B1(new_n897_), .B2(new_n904_), .ZN(new_n905_));
  AND2_X1   g544(.A1(new_n903_), .A2(G8), .ZN(new_n906_));
  AOI21_X1  g545(.A(new_n902_), .B1(new_n906_), .B2(new_n898_), .ZN(new_n907_));
  OAI21_X1  g546(.A(KEYINPUT61), .B1(new_n907_), .B2(new_n904_), .ZN(new_n908_));
  INV_X1    g547(.A(KEYINPUT54), .ZN(new_n909_));
  NAND3_X1  g548(.A1(new_n888_), .A2(new_n909_), .A3(new_n612_), .ZN(new_n910_));
  INV_X1    g549(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g550(.A1(new_n888_), .A2(G2078), .ZN(new_n912_));
  NOR2_X1   g551(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g552(.A(new_n909_), .B1(new_n888_), .B2(new_n612_), .ZN(new_n914_));
  INV_X1    g553(.A(new_n914_), .ZN(new_n915_));
  AOI21_X1  g554(.A(G301), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g555(.A1(new_n898_), .A2(G8), .A3(new_n903_), .ZN(new_n917_));
  NAND3_X1  g556(.A1(new_n917_), .A2(new_n899_), .A3(new_n901_), .ZN(new_n918_));
  NAND3_X1  g557(.A1(new_n906_), .A2(new_n902_), .A3(new_n898_), .ZN(new_n919_));
  INV_X1    g558(.A(KEYINPUT61), .ZN(new_n920_));
  NAND3_X1  g559(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  NAND4_X1  g560(.A1(new_n897_), .A2(new_n908_), .A3(new_n916_), .A4(new_n921_), .ZN(new_n922_));
  OR2_X1    g561(.A1(new_n896_), .A2(KEYINPUT62), .ZN(new_n923_));
  INV_X1    g562(.A(new_n892_), .ZN(new_n924_));
  NAND2_X1  g563(.A1(new_n896_), .A2(KEYINPUT62), .ZN(new_n925_));
  NAND3_X1  g564(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  NAND3_X1  g565(.A1(new_n905_), .A2(new_n922_), .A3(new_n926_), .ZN(new_n927_));
  NAND3_X1  g566(.A1(new_n835_), .A2(G2067), .A3(new_n882_), .ZN(new_n928_));
  NAND2_X1  g567(.A1(new_n888_), .A2(G1348), .ZN(new_n929_));
  NAND3_X1  g568(.A1(new_n928_), .A2(new_n929_), .A3(new_n520_), .ZN(new_n930_));
  NAND2_X1  g569(.A1(new_n930_), .A2(KEYINPUT56), .ZN(new_n931_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n932_));
  NAND4_X1  g571(.A1(new_n928_), .A2(new_n929_), .A3(new_n932_), .A4(new_n520_), .ZN(new_n933_));
  NAND2_X1  g572(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g573(.A1(new_n835_), .A2(G2072), .A3(new_n882_), .ZN(new_n935_));
  NAND2_X1  g574(.A1(new_n888_), .A2(G1956), .ZN(new_n936_));
  AND3_X1   g575(.A1(new_n935_), .A2(new_n936_), .A3(new_n487_), .ZN(new_n937_));
  AOI21_X1  g576(.A(new_n487_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n938_));
  NOR2_X1   g577(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g578(.A1(new_n934_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g579(.A1(new_n940_), .A2(KEYINPUT57), .ZN(new_n941_));
  XOR2_X1   g580(.A(new_n937_), .B(KEYINPUT58), .Z(new_n942_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n943_));
  NAND3_X1  g582(.A1(new_n934_), .A2(new_n939_), .A3(new_n943_), .ZN(new_n944_));
  XOR2_X1   g583(.A(KEYINPUT59), .B(G1341), .Z(new_n945_));
  NAND2_X1  g584(.A1(new_n888_), .A2(new_n945_), .ZN(new_n946_));
  OR2_X1    g585(.A1(new_n946_), .A2(KEYINPUT60), .ZN(new_n947_));
  NAND2_X1  g586(.A1(new_n946_), .A2(KEYINPUT60), .ZN(new_n948_));
  OAI211_X1 g587(.A(new_n947_), .B(new_n948_), .C1(G1996), .C2(new_n888_), .ZN(new_n949_));
  NAND2_X1  g588(.A1(new_n928_), .A2(new_n929_), .ZN(new_n950_));
  AOI21_X1  g589(.A(new_n474_), .B1(new_n950_), .B2(new_n530_), .ZN(new_n951_));
  NAND4_X1  g590(.A1(new_n949_), .A2(new_n939_), .A3(new_n930_), .A4(new_n951_), .ZN(new_n952_));
  NAND4_X1  g591(.A1(new_n941_), .A2(new_n942_), .A3(new_n944_), .A4(new_n952_), .ZN(new_n953_));
  NOR2_X1   g592(.A1(new_n907_), .A2(new_n904_), .ZN(new_n954_));
  NAND2_X1  g593(.A1(new_n897_), .A2(new_n954_), .ZN(new_n955_));
  INV_X1    g594(.A(new_n912_), .ZN(new_n956_));
  NAND2_X1  g595(.A1(new_n956_), .A2(new_n910_), .ZN(new_n957_));
  OAI21_X1  g596(.A(new_n609_), .B1(new_n957_), .B2(new_n914_), .ZN(new_n958_));
  NAND4_X1  g597(.A1(new_n915_), .A2(new_n956_), .A3(G301), .A4(new_n910_), .ZN(new_n959_));
  NAND2_X1  g598(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n961_));
  NAND2_X1  g600(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  NAND3_X1  g601(.A1(new_n958_), .A2(KEYINPUT55), .A3(new_n959_), .ZN(new_n963_));
  AOI21_X1  g602(.A(new_n955_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  AOI21_X1  g603(.A(new_n927_), .B1(new_n953_), .B2(new_n964_), .ZN(new_n965_));
  OR2_X1    g604(.A1(new_n851_), .A2(new_n854_), .ZN(new_n966_));
  NAND4_X1  g605(.A1(new_n966_), .A2(new_n855_), .A3(new_n859_), .A4(new_n862_), .ZN(new_n967_));
  OAI21_X1  g606(.A(new_n868_), .B1(new_n965_), .B2(new_n967_), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g607(.A1(new_n595_), .A2(new_n596_), .A3(G319), .ZN(new_n970_));
  NOR2_X1   g608(.A1(new_n970_), .A2(G401), .ZN(new_n971_));
  NAND2_X1  g609(.A1(new_n971_), .A2(new_n826_), .ZN(new_n972_));
  NAND2_X1  g610(.A1(new_n782_), .A2(new_n788_), .ZN(new_n973_));
  NAND2_X1  g611(.A1(new_n973_), .A2(new_n734_), .ZN(new_n974_));
  INV_X1    g612(.A(G227), .ZN(new_n975_));
  NAND3_X1  g613(.A1(new_n974_), .A2(KEYINPUT63), .A3(new_n975_), .ZN(new_n976_));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n977_));
  OAI21_X1  g615(.A(new_n977_), .B1(G395), .B2(G227), .ZN(new_n978_));
  AOI21_X1  g616(.A(new_n972_), .B1(new_n976_), .B2(new_n978_), .ZN(G308));
  AND2_X1   g617(.A1(new_n971_), .A2(new_n826_), .ZN(new_n980_));
  AOI21_X1  g618(.A(KEYINPUT63), .B1(new_n974_), .B2(new_n975_), .ZN(new_n981_));
  NOR3_X1   g619(.A1(G395), .A2(new_n977_), .A3(G227), .ZN(new_n982_));
  OAI21_X1  g620(.A(new_n980_), .B1(new_n981_), .B2(new_n982_), .ZN(G225));
endmodule


