//Secret key is'0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_c1908" written by ABC on Wed Oct 26 13:45:21 2022

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110,
    G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146,
    G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478,
    G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104,
    G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140,
    G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472,
    G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n574_, new_n575_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_;
  INV_X1    g000(.A(G472), .ZN(new_n123_));
  INV_X1    g001(.A(G953), .ZN(new_n124_));
  NAND2_X1  g002(.A1(new_n124_), .A2(KEYINPUT10), .ZN(new_n125_));
  INV_X1    g003(.A(KEYINPUT10), .ZN(new_n126_));
  NAND2_X1  g004(.A1(new_n126_), .A2(G953), .ZN(new_n127_));
  NAND2_X1  g005(.A1(new_n125_), .A2(new_n127_), .ZN(new_n128_));
  INV_X1    g006(.A(G237), .ZN(new_n129_));
  NAND2_X1  g007(.A1(new_n129_), .A2(G210), .ZN(new_n130_));
  OAI21_X1  g008(.A(KEYINPUT28), .B1(new_n128_), .B2(new_n130_), .ZN(new_n131_));
  INV_X1    g009(.A(new_n131_), .ZN(new_n132_));
  NOR3_X1   g010(.A1(new_n128_), .A2(KEYINPUT28), .A3(new_n130_), .ZN(new_n133_));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G101), .ZN(new_n134_));
  INV_X1    g012(.A(new_n134_), .ZN(new_n135_));
  NOR3_X1   g013(.A1(new_n132_), .A2(new_n133_), .A3(new_n135_), .ZN(new_n136_));
  INV_X1    g014(.A(new_n133_), .ZN(new_n137_));
  AOI21_X1  g015(.A(new_n134_), .B1(new_n137_), .B2(new_n131_), .ZN(new_n138_));
  NOR2_X1   g016(.A1(new_n136_), .A2(new_n138_), .ZN(new_n139_));
  INV_X1    g017(.A(G143), .ZN(new_n140_));
  INV_X1    g018(.A(G146), .ZN(new_n141_));
  NAND2_X1  g019(.A1(new_n140_), .A2(new_n141_), .ZN(new_n142_));
  NAND2_X1  g020(.A1(G143), .A2(G146), .ZN(new_n143_));
  NAND3_X1  g021(.A1(new_n142_), .A2(G128), .A3(new_n143_), .ZN(new_n144_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n145_));
  NAND2_X1  g023(.A1(new_n144_), .A2(new_n145_), .ZN(new_n146_));
  NAND4_X1  g024(.A1(new_n142_), .A2(KEYINPUT3), .A3(G128), .A4(new_n143_), .ZN(new_n147_));
  AND2_X1   g025(.A1(new_n146_), .A2(new_n147_), .ZN(new_n148_));
  XNOR2_X1  g026(.A(G134), .B(G137), .ZN(new_n149_));
  INV_X1    g027(.A(G131), .ZN(new_n150_));
  XNOR2_X1  g028(.A(new_n149_), .B(new_n150_), .ZN(new_n151_));
  INV_X1    g029(.A(G128), .ZN(new_n152_));
  AND2_X1   g030(.A1(G143), .A2(G146), .ZN(new_n153_));
  NOR2_X1   g031(.A1(G143), .A2(G146), .ZN(new_n154_));
  OAI21_X1  g032(.A(new_n152_), .B1(new_n153_), .B2(new_n154_), .ZN(new_n155_));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n156_));
  NAND2_X1  g034(.A1(new_n155_), .A2(new_n156_), .ZN(new_n157_));
  OAI211_X1 g035(.A(KEYINPUT2), .B(new_n152_), .C1(new_n153_), .C2(new_n154_), .ZN(new_n158_));
  NAND2_X1  g036(.A1(new_n157_), .A2(new_n158_), .ZN(new_n159_));
  NAND3_X1  g037(.A1(new_n148_), .A2(new_n151_), .A3(new_n159_), .ZN(new_n160_));
  NOR2_X1   g038(.A1(G116), .A2(G119), .ZN(new_n161_));
  INV_X1    g039(.A(new_n161_), .ZN(new_n162_));
  NAND2_X1  g040(.A1(G116), .A2(G119), .ZN(new_n163_));
  NAND3_X1  g041(.A1(new_n162_), .A2(G113), .A3(new_n163_), .ZN(new_n164_));
  INV_X1    g042(.A(G113), .ZN(new_n165_));
  INV_X1    g043(.A(new_n163_), .ZN(new_n166_));
  OAI21_X1  g044(.A(new_n165_), .B1(new_n166_), .B2(new_n161_), .ZN(new_n167_));
  NAND2_X1  g045(.A1(new_n164_), .A2(new_n167_), .ZN(new_n168_));
  XNOR2_X1  g046(.A(new_n149_), .B(G131), .ZN(new_n169_));
  NAND2_X1  g047(.A1(new_n155_), .A2(new_n144_), .ZN(new_n170_));
  NAND2_X1  g048(.A1(new_n169_), .A2(new_n170_), .ZN(new_n171_));
  NAND3_X1  g049(.A1(new_n160_), .A2(new_n168_), .A3(new_n171_), .ZN(new_n172_));
  INV_X1    g050(.A(new_n172_), .ZN(new_n173_));
  AOI21_X1  g051(.A(new_n168_), .B1(new_n160_), .B2(new_n171_), .ZN(new_n174_));
  OAI21_X1  g052(.A(new_n139_), .B1(new_n173_), .B2(new_n174_), .ZN(new_n175_));
  NAND2_X1  g053(.A1(new_n160_), .A2(new_n171_), .ZN(new_n176_));
  INV_X1    g054(.A(new_n168_), .ZN(new_n177_));
  NAND2_X1  g055(.A1(new_n176_), .A2(new_n177_), .ZN(new_n178_));
  OR2_X1    g056(.A1(new_n136_), .A2(new_n138_), .ZN(new_n179_));
  NAND3_X1  g057(.A1(new_n178_), .A2(new_n172_), .A3(new_n179_), .ZN(new_n180_));
  NAND2_X1  g058(.A1(new_n175_), .A2(new_n180_), .ZN(new_n181_));
  INV_X1    g059(.A(G902), .ZN(new_n182_));
  AOI21_X1  g060(.A(new_n123_), .B1(new_n181_), .B2(new_n182_), .ZN(new_n183_));
  AOI211_X1 g061(.A(G472), .B(G902), .C1(new_n175_), .C2(new_n180_), .ZN(new_n184_));
  NOR2_X1   g062(.A1(new_n183_), .A2(new_n184_), .ZN(new_n185_));
  AND2_X1   g063(.A1(new_n125_), .A2(new_n127_), .ZN(new_n186_));
  NAND4_X1  g064(.A1(new_n186_), .A2(G137), .A3(G221), .A4(G234), .ZN(new_n187_));
  INV_X1    g065(.A(G137), .ZN(new_n188_));
  NAND2_X1  g066(.A1(G221), .A2(G234), .ZN(new_n189_));
  OAI21_X1  g067(.A(new_n188_), .B1(new_n128_), .B2(new_n189_), .ZN(new_n190_));
  NAND2_X1  g068(.A1(new_n187_), .A2(new_n190_), .ZN(new_n191_));
  INV_X1    g069(.A(new_n191_), .ZN(new_n192_));
  NAND2_X1  g070(.A1(G125), .A2(G140), .ZN(new_n193_));
  NOR2_X1   g071(.A1(G125), .A2(G140), .ZN(new_n194_));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n195_));
  OAI21_X1  g073(.A(new_n193_), .B1(new_n194_), .B2(new_n195_), .ZN(new_n196_));
  INV_X1    g074(.A(new_n193_), .ZN(new_n197_));
  NAND2_X1  g075(.A1(new_n197_), .A2(KEYINPUT23), .ZN(new_n198_));
  NAND2_X1  g076(.A1(new_n196_), .A2(new_n198_), .ZN(new_n199_));
  NAND2_X1  g077(.A1(new_n199_), .A2(new_n141_), .ZN(new_n200_));
  OR2_X1    g078(.A1(G119), .A2(G128), .ZN(new_n201_));
  NAND2_X1  g079(.A1(G119), .A2(G128), .ZN(new_n202_));
  NAND2_X1  g080(.A1(new_n201_), .A2(new_n202_), .ZN(new_n203_));
  INV_X1    g081(.A(G110), .ZN(new_n204_));
  NAND2_X1  g082(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g083(.A1(new_n201_), .A2(G110), .A3(new_n202_), .ZN(new_n206_));
  NAND2_X1  g084(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g085(.A(KEYINPUT21), .B1(new_n197_), .B2(new_n194_), .ZN(new_n208_));
  INV_X1    g086(.A(G140), .ZN(new_n209_));
  NOR3_X1   g087(.A1(new_n209_), .A2(KEYINPUT21), .A3(G125), .ZN(new_n210_));
  INV_X1    g088(.A(new_n210_), .ZN(new_n211_));
  NAND3_X1  g089(.A1(new_n208_), .A2(new_n211_), .A3(G146), .ZN(new_n212_));
  NAND3_X1  g090(.A1(new_n200_), .A2(new_n207_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g091(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n215_));
  INV_X1    g093(.A(G125), .ZN(new_n216_));
  NAND2_X1  g094(.A1(new_n216_), .A2(new_n209_), .ZN(new_n217_));
  AOI21_X1  g095(.A(new_n215_), .B1(new_n217_), .B2(new_n193_), .ZN(new_n218_));
  OAI21_X1  g096(.A(new_n141_), .B1(new_n218_), .B2(new_n210_), .ZN(new_n219_));
  AOI21_X1  g097(.A(new_n207_), .B1(new_n212_), .B2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g098(.A(new_n192_), .B1(new_n214_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g099(.A1(new_n219_), .A2(new_n212_), .ZN(new_n222_));
  NAND3_X1  g100(.A1(new_n222_), .A2(new_n206_), .A3(new_n205_), .ZN(new_n223_));
  NAND3_X1  g101(.A1(new_n223_), .A2(new_n191_), .A3(new_n213_), .ZN(new_n224_));
  NAND3_X1  g102(.A1(new_n221_), .A2(new_n224_), .A3(new_n182_), .ZN(new_n225_));
  INV_X1    g103(.A(G217), .ZN(new_n226_));
  AOI21_X1  g104(.A(new_n226_), .B1(G234), .B2(new_n182_), .ZN(new_n227_));
  NAND2_X1  g105(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g106(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n229_));
  INV_X1    g107(.A(KEYINPUT26), .ZN(new_n230_));
  NAND3_X1  g108(.A1(new_n225_), .A2(new_n230_), .A3(new_n227_), .ZN(new_n231_));
  INV_X1    g109(.A(new_n227_), .ZN(new_n232_));
  NAND3_X1  g110(.A1(new_n221_), .A2(new_n224_), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g111(.A1(new_n233_), .A2(G902), .ZN(new_n234_));
  NAND3_X1  g112(.A1(new_n229_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n235_));
  NOR2_X1   g113(.A1(new_n185_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g114(.A(G113), .B(G122), .ZN(new_n237_));
  XNOR2_X1  g115(.A(new_n237_), .B(G104), .ZN(new_n238_));
  NAND3_X1  g116(.A1(new_n217_), .A2(G146), .A3(new_n193_), .ZN(new_n239_));
  NAND2_X1  g117(.A1(new_n200_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g118(.A1(new_n129_), .A2(new_n124_), .A3(G214), .ZN(new_n241_));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n242_));
  AOI21_X1  g120(.A(G143), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g121(.A(G214), .ZN(new_n244_));
  NOR3_X1   g122(.A1(new_n244_), .A2(G237), .A3(G953), .ZN(new_n245_));
  NAND2_X1  g123(.A1(new_n245_), .A2(KEYINPUT22), .ZN(new_n246_));
  NAND2_X1  g124(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g125(.A1(new_n244_), .A2(G237), .ZN(new_n248_));
  NAND4_X1  g126(.A1(new_n248_), .A2(new_n125_), .A3(new_n127_), .A4(G143), .ZN(new_n249_));
  NAND3_X1  g127(.A1(new_n247_), .A2(new_n150_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g128(.A(new_n249_), .B1(G143), .B2(new_n245_), .ZN(new_n251_));
  NAND2_X1  g129(.A1(new_n251_), .A2(G131), .ZN(new_n252_));
  NAND3_X1  g130(.A1(new_n240_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g131(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g132(.A1(new_n200_), .A2(new_n212_), .ZN(new_n255_));
  NAND3_X1  g133(.A1(new_n248_), .A2(new_n125_), .A3(new_n127_), .ZN(new_n256_));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n257_));
  OAI21_X1  g135(.A(new_n256_), .B1(new_n257_), .B2(G143), .ZN(new_n258_));
  NOR2_X1   g136(.A1(new_n257_), .A2(G143), .ZN(new_n259_));
  NAND4_X1  g137(.A1(new_n248_), .A2(new_n259_), .A3(new_n125_), .A4(new_n127_), .ZN(new_n260_));
  NAND3_X1  g138(.A1(new_n258_), .A2(G131), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g139(.A(new_n255_), .B1(new_n250_), .B2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g140(.A(new_n238_), .B1(new_n254_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g141(.A1(new_n263_), .A2(KEYINPUT25), .ZN(new_n264_));
  INV_X1    g142(.A(new_n238_), .ZN(new_n265_));
  NAND2_X1  g143(.A1(new_n250_), .A2(new_n261_), .ZN(new_n266_));
  INV_X1    g144(.A(new_n255_), .ZN(new_n267_));
  NAND2_X1  g145(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g146(.A(new_n265_), .B1(new_n268_), .B2(new_n253_), .ZN(new_n269_));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n270_));
  NAND2_X1  g148(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g149(.A1(new_n256_), .A2(new_n140_), .ZN(new_n272_));
  NAND2_X1  g150(.A1(new_n272_), .A2(new_n249_), .ZN(new_n273_));
  NAND2_X1  g151(.A1(new_n273_), .A2(G131), .ZN(new_n274_));
  NAND2_X1  g152(.A1(new_n274_), .A2(new_n250_), .ZN(new_n275_));
  AND2_X1   g153(.A1(new_n219_), .A2(new_n212_), .ZN(new_n276_));
  NAND2_X1  g154(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g155(.A1(new_n277_), .A2(new_n265_), .A3(new_n253_), .ZN(new_n278_));
  NAND3_X1  g156(.A1(new_n264_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n279_));
  NOR2_X1   g157(.A1(G475), .A2(G902), .ZN(new_n280_));
  AOI21_X1  g158(.A(new_n222_), .B1(new_n274_), .B2(new_n250_), .ZN(new_n281_));
  NOR3_X1   g159(.A1(new_n254_), .A2(new_n281_), .A3(new_n238_), .ZN(new_n282_));
  AOI21_X1  g160(.A(new_n265_), .B1(new_n277_), .B2(new_n253_), .ZN(new_n283_));
  OAI21_X1  g161(.A(new_n182_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  AOI22_X1  g162(.A1(new_n279_), .A2(new_n280_), .B1(new_n284_), .B2(G475), .ZN(new_n285_));
  XNOR2_X1  g163(.A(G128), .B(G143), .ZN(new_n286_));
  INV_X1    g164(.A(G134), .ZN(new_n287_));
  NAND2_X1  g165(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g166(.A1(G116), .A2(G122), .ZN(new_n289_));
  NAND2_X1  g167(.A1(G116), .A2(G122), .ZN(new_n290_));
  AOI21_X1  g168(.A(G107), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g169(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g170(.A1(new_n289_), .A2(G107), .A3(new_n290_), .ZN(new_n293_));
  NAND2_X1  g171(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g172(.A(KEYINPUT17), .ZN(new_n295_));
  NAND2_X1  g173(.A1(new_n286_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g174(.A1(new_n152_), .A2(G143), .ZN(new_n297_));
  AOI21_X1  g175(.A(new_n287_), .B1(new_n297_), .B2(KEYINPUT17), .ZN(new_n298_));
  AND3_X1   g176(.A1(new_n296_), .A2(KEYINPUT18), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g177(.A(KEYINPUT18), .B1(new_n296_), .B2(new_n298_), .ZN(new_n300_));
  OAI211_X1 g178(.A(new_n288_), .B(new_n294_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g179(.A(KEYINPUT19), .B1(new_n286_), .B2(new_n287_), .ZN(new_n302_));
  OAI21_X1  g180(.A(new_n302_), .B1(new_n287_), .B2(new_n286_), .ZN(new_n303_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n304_));
  OAI21_X1  g182(.A(new_n293_), .B1(new_n291_), .B2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g183(.A1(new_n289_), .A2(KEYINPUT20), .A3(G107), .A4(new_n290_), .ZN(new_n306_));
  INV_X1    g184(.A(new_n286_), .ZN(new_n307_));
  NAND3_X1  g185(.A1(new_n307_), .A2(KEYINPUT19), .A3(G134), .ZN(new_n308_));
  NAND4_X1  g186(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g187(.A(G234), .ZN(new_n310_));
  NOR3_X1   g188(.A1(new_n226_), .A2(new_n310_), .A3(G953), .ZN(new_n311_));
  AND3_X1   g189(.A1(new_n301_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g190(.A(new_n311_), .B1(new_n301_), .B2(new_n309_), .ZN(new_n313_));
  OAI21_X1  g191(.A(new_n182_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g192(.A1(new_n314_), .A2(G478), .ZN(new_n315_));
  INV_X1    g193(.A(G478), .ZN(new_n316_));
  OAI211_X1 g194(.A(new_n316_), .B(new_n182_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n317_));
  NAND2_X1  g195(.A1(G234), .A2(G237), .ZN(new_n318_));
  NAND3_X1  g196(.A1(new_n186_), .A2(G952), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g197(.A(new_n182_), .B1(G234), .B2(G237), .ZN(new_n320_));
  INV_X1    g198(.A(G898), .ZN(new_n321_));
  NAND3_X1  g199(.A1(new_n320_), .A2(new_n321_), .A3(G953), .ZN(new_n322_));
  NAND2_X1  g200(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  AND4_X1   g201(.A1(new_n285_), .A2(new_n315_), .A3(new_n317_), .A4(new_n323_), .ZN(new_n324_));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325_));
  XNOR2_X1  g203(.A(new_n325_), .B(KEYINPUT0), .ZN(new_n326_));
  OAI21_X1  g204(.A(G210), .B1(G237), .B2(G902), .ZN(new_n327_));
  XNOR2_X1  g205(.A(new_n327_), .B(KEYINPUT9), .ZN(new_n328_));
  NAND2_X1  g206(.A1(new_n124_), .A2(G224), .ZN(new_n329_));
  XNOR2_X1  g207(.A(new_n329_), .B(KEYINPUT1), .ZN(new_n330_));
  INV_X1    g208(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g209(.A1(new_n170_), .A2(G125), .ZN(new_n332_));
  NAND3_X1  g210(.A1(new_n159_), .A2(new_n146_), .A3(new_n147_), .ZN(new_n333_));
  AOI21_X1  g211(.A(new_n332_), .B1(new_n333_), .B2(G125), .ZN(new_n334_));
  OAI21_X1  g212(.A(new_n331_), .B1(new_n334_), .B2(KEYINPUT6), .ZN(new_n335_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n336_));
  AOI21_X1  g214(.A(new_n216_), .B1(new_n148_), .B2(new_n159_), .ZN(new_n337_));
  OAI211_X1 g215(.A(new_n336_), .B(new_n330_), .C1(new_n337_), .C2(new_n332_), .ZN(new_n338_));
  INV_X1    g216(.A(G101), .ZN(new_n339_));
  AND2_X1   g217(.A1(G104), .A2(G107), .ZN(new_n340_));
  NOR2_X1   g218(.A1(G104), .A2(G107), .ZN(new_n341_));
  OAI21_X1  g219(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g220(.A(G104), .ZN(new_n343_));
  INV_X1    g221(.A(G107), .ZN(new_n344_));
  NAND2_X1  g222(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g223(.A1(G104), .A2(G107), .ZN(new_n346_));
  NAND3_X1  g224(.A1(new_n345_), .A2(G101), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g225(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g226(.A1(new_n164_), .A2(new_n167_), .A3(KEYINPUT5), .ZN(new_n349_));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n350_));
  NAND4_X1  g228(.A1(new_n162_), .A2(new_n350_), .A3(G113), .A4(new_n163_), .ZN(new_n351_));
  AOI21_X1  g229(.A(new_n348_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g230(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n354_));
  NAND2_X1  g232(.A1(new_n168_), .A2(new_n348_), .ZN(new_n355_));
  NAND3_X1  g233(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g234(.A1(new_n335_), .A2(new_n338_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g235(.A1(new_n349_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n358_));
  OAI21_X1  g236(.A(new_n358_), .B1(new_n352_), .B2(KEYINPUT7), .ZN(new_n359_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n360_));
  NAND4_X1  g238(.A1(new_n349_), .A2(new_n360_), .A3(new_n348_), .A4(new_n351_), .ZN(new_n361_));
  NAND2_X1  g239(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g240(.A(new_n354_), .ZN(new_n363_));
  NAND2_X1  g241(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g242(.A(KEYINPUT8), .ZN(new_n365_));
  NAND2_X1  g243(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g244(.A1(new_n362_), .A2(KEYINPUT8), .A3(new_n363_), .ZN(new_n367_));
  AOI21_X1  g245(.A(new_n357_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g246(.A(new_n355_), .ZN(new_n369_));
  OAI21_X1  g247(.A(new_n363_), .B1(new_n352_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g248(.A1(new_n356_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n372_));
  NAND2_X1  g250(.A1(new_n331_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g251(.A1(new_n330_), .A2(KEYINPUT4), .ZN(new_n374_));
  NAND3_X1  g252(.A1(new_n334_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  OAI211_X1 g253(.A(new_n372_), .B(new_n331_), .C1(new_n337_), .C2(new_n332_), .ZN(new_n376_));
  NAND3_X1  g254(.A1(new_n371_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g255(.A1(new_n377_), .A2(new_n182_), .ZN(new_n378_));
  OAI21_X1  g256(.A(new_n328_), .B1(new_n368_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g257(.A(new_n356_), .ZN(new_n380_));
  OAI21_X1  g258(.A(new_n336_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n381_));
  AOI21_X1  g259(.A(new_n380_), .B1(new_n381_), .B2(new_n331_), .ZN(new_n382_));
  AOI21_X1  g260(.A(KEYINPUT8), .B1(new_n362_), .B2(new_n363_), .ZN(new_n383_));
  AOI211_X1 g261(.A(new_n365_), .B(new_n354_), .C1(new_n359_), .C2(new_n361_), .ZN(new_n384_));
  OAI211_X1 g262(.A(new_n382_), .B(new_n338_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  INV_X1    g263(.A(new_n378_), .ZN(new_n386_));
  INV_X1    g264(.A(new_n328_), .ZN(new_n387_));
  NAND3_X1  g265(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g266(.A(new_n326_), .B1(new_n379_), .B2(new_n388_), .ZN(new_n389_));
  AND2_X1   g267(.A1(new_n324_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g268(.A1(new_n142_), .A2(new_n143_), .ZN(new_n391_));
  AOI21_X1  g269(.A(KEYINPUT2), .B1(new_n391_), .B2(new_n152_), .ZN(new_n392_));
  INV_X1    g270(.A(new_n158_), .ZN(new_n393_));
  NOR2_X1   g271(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g272(.A1(new_n146_), .A2(new_n147_), .ZN(new_n395_));
  OAI21_X1  g273(.A(new_n348_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g274(.A1(new_n155_), .A2(new_n144_), .A3(new_n342_), .A4(new_n347_), .ZN(new_n397_));
  INV_X1    g275(.A(KEYINPUT11), .ZN(new_n398_));
  NAND2_X1  g276(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g277(.A(new_n170_), .ZN(new_n400_));
  AND2_X1   g278(.A1(new_n342_), .A2(new_n347_), .ZN(new_n401_));
  NAND3_X1  g279(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT11), .ZN(new_n402_));
  NAND4_X1  g280(.A1(new_n396_), .A2(new_n169_), .A3(new_n399_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g281(.A1(new_n403_), .A2(KEYINPUT12), .ZN(new_n404_));
  NAND2_X1  g282(.A1(new_n402_), .A2(new_n399_), .ZN(new_n405_));
  INV_X1    g283(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n407_));
  NAND4_X1  g285(.A1(new_n406_), .A2(new_n407_), .A3(new_n169_), .A4(new_n396_), .ZN(new_n408_));
  INV_X1    g286(.A(new_n396_), .ZN(new_n409_));
  OAI21_X1  g287(.A(new_n151_), .B1(new_n409_), .B2(new_n405_), .ZN(new_n410_));
  NAND3_X1  g288(.A1(new_n404_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g289(.A1(new_n186_), .A2(G227), .ZN(new_n412_));
  XNOR2_X1  g290(.A(G110), .B(G140), .ZN(new_n413_));
  XNOR2_X1  g291(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g292(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g293(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  AOI22_X1  g294(.A1(new_n155_), .A2(new_n144_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n417_));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n418_));
  AOI21_X1  g296(.A(new_n417_), .B1(new_n418_), .B2(new_n397_), .ZN(new_n419_));
  NAND3_X1  g297(.A1(new_n170_), .A2(new_n348_), .A3(new_n418_), .ZN(new_n420_));
  INV_X1    g298(.A(new_n420_), .ZN(new_n421_));
  OAI21_X1  g299(.A(new_n151_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n423_));
  NAND2_X1  g301(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g302(.A1(new_n397_), .A2(new_n418_), .ZN(new_n425_));
  NAND2_X1  g303(.A1(new_n170_), .A2(new_n348_), .ZN(new_n426_));
  NAND2_X1  g304(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g305(.A1(new_n427_), .A2(new_n420_), .ZN(new_n428_));
  NAND3_X1  g306(.A1(new_n428_), .A2(KEYINPUT14), .A3(new_n151_), .ZN(new_n429_));
  NAND2_X1  g307(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  AND2_X1   g308(.A1(new_n403_), .A2(new_n414_), .ZN(new_n431_));
  NAND2_X1  g309(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g310(.A1(new_n416_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g311(.A(G469), .ZN(new_n434_));
  NAND3_X1  g312(.A1(new_n433_), .A2(new_n434_), .A3(new_n182_), .ZN(new_n435_));
  AOI21_X1  g313(.A(new_n414_), .B1(new_n430_), .B2(new_n403_), .ZN(new_n436_));
  AND4_X1   g314(.A1(new_n414_), .A2(new_n404_), .A3(new_n408_), .A4(new_n410_), .ZN(new_n437_));
  OAI211_X1 g315(.A(KEYINPUT15), .B(new_n182_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g316(.A1(new_n438_), .A2(G469), .ZN(new_n439_));
  AOI21_X1  g317(.A(KEYINPUT14), .B1(new_n428_), .B2(new_n151_), .ZN(new_n440_));
  AOI211_X1 g318(.A(new_n423_), .B(new_n169_), .C1(new_n427_), .C2(new_n420_), .ZN(new_n441_));
  OAI21_X1  g319(.A(new_n403_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g320(.A1(new_n442_), .A2(new_n415_), .ZN(new_n443_));
  NAND4_X1  g321(.A1(new_n404_), .A2(new_n408_), .A3(new_n410_), .A4(new_n414_), .ZN(new_n444_));
  NAND2_X1  g322(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g323(.A(KEYINPUT15), .B1(new_n445_), .B2(new_n182_), .ZN(new_n446_));
  OAI21_X1  g324(.A(new_n435_), .B1(new_n439_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g325(.A(G221), .B1(new_n310_), .B2(G902), .ZN(new_n448_));
  AND3_X1   g326(.A1(new_n447_), .A2(KEYINPUT16), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g327(.A(KEYINPUT16), .B1(new_n447_), .B2(new_n448_), .ZN(new_n450_));
  OAI211_X1 g328(.A(new_n236_), .B(new_n390_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g329(.A1(new_n451_), .A2(KEYINPUT29), .ZN(new_n452_));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n453_));
  AOI22_X1  g331(.A1(new_n411_), .A2(new_n415_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n454_));
  NOR3_X1   g332(.A1(new_n454_), .A2(G469), .A3(G902), .ZN(new_n455_));
  AOI21_X1  g333(.A(G902), .B1(new_n443_), .B2(new_n444_), .ZN(new_n456_));
  AOI21_X1  g334(.A(new_n434_), .B1(new_n456_), .B2(KEYINPUT15), .ZN(new_n457_));
  OAI21_X1  g335(.A(new_n182_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n458_));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n459_));
  NAND2_X1  g337(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g338(.A(new_n455_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g339(.A(new_n448_), .ZN(new_n462_));
  OAI21_X1  g340(.A(new_n453_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g341(.A1(new_n447_), .A2(KEYINPUT16), .A3(new_n448_), .ZN(new_n464_));
  NAND2_X1  g342(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n466_));
  NAND4_X1  g344(.A1(new_n465_), .A2(new_n466_), .A3(new_n236_), .A4(new_n390_), .ZN(new_n467_));
  NAND2_X1  g345(.A1(new_n452_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g346(.A(new_n468_), .B(G101), .ZN(G3));
  NOR2_X1   g347(.A1(new_n449_), .A2(new_n450_), .ZN(new_n470_));
  NOR3_X1   g348(.A1(new_n235_), .A2(new_n183_), .A3(new_n184_), .ZN(new_n471_));
  INV_X1    g349(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g350(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g351(.A1(new_n379_), .A2(new_n388_), .ZN(new_n474_));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n475_));
  NAND2_X1  g353(.A1(new_n317_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g354(.A1(new_n301_), .A2(new_n309_), .ZN(new_n477_));
  INV_X1    g355(.A(new_n311_), .ZN(new_n478_));
  NAND2_X1  g356(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g357(.A1(new_n301_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n480_));
  NAND2_X1  g358(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g359(.A1(new_n481_), .A2(KEYINPUT30), .A3(new_n316_), .A4(new_n182_), .ZN(new_n482_));
  NAND3_X1  g360(.A1(new_n476_), .A2(new_n482_), .A3(new_n315_), .ZN(new_n483_));
  NOR2_X1   g361(.A1(new_n285_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g362(.A(new_n326_), .ZN(new_n485_));
  NAND4_X1  g363(.A1(new_n474_), .A2(new_n484_), .A3(new_n485_), .A4(new_n323_), .ZN(new_n486_));
  INV_X1    g364(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g365(.A1(new_n473_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g366(.A(new_n488_), .B(G104), .ZN(G6));
  NOR3_X1   g367(.A1(new_n368_), .A2(new_n328_), .A3(new_n378_), .ZN(new_n490_));
  AOI21_X1  g368(.A(new_n387_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n491_));
  OAI211_X1 g369(.A(new_n485_), .B(new_n323_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g370(.A(G475), .ZN(new_n493_));
  OAI21_X1  g371(.A(new_n238_), .B1(new_n254_), .B2(new_n281_), .ZN(new_n494_));
  AOI21_X1  g372(.A(G902), .B1(new_n494_), .B2(new_n278_), .ZN(new_n495_));
  AOI21_X1  g373(.A(new_n493_), .B1(new_n495_), .B2(KEYINPUT31), .ZN(new_n496_));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n497_));
  NAND2_X1  g375(.A1(new_n284_), .A2(new_n497_), .ZN(new_n498_));
  AOI22_X1  g376(.A1(new_n496_), .A2(new_n498_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n499_));
  NAND2_X1  g377(.A1(new_n315_), .A2(new_n317_), .ZN(new_n500_));
  NAND2_X1  g378(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g379(.A1(new_n492_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g380(.A1(new_n473_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G107), .Z(new_n504_));
  XNOR2_X1  g382(.A(new_n503_), .B(new_n504_), .ZN(G9));
  NAND2_X1  g383(.A1(new_n233_), .A2(KEYINPUT33), .ZN(new_n506_));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n507_));
  NAND4_X1  g385(.A1(new_n221_), .A2(new_n224_), .A3(new_n507_), .A4(new_n232_), .ZN(new_n508_));
  NAND3_X1  g386(.A1(new_n506_), .A2(new_n182_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g387(.A1(new_n509_), .A2(new_n228_), .ZN(new_n510_));
  AOI21_X1  g388(.A(KEYINPUT34), .B1(new_n185_), .B2(new_n510_), .ZN(new_n511_));
  NOR3_X1   g389(.A1(new_n173_), .A2(new_n174_), .A3(new_n139_), .ZN(new_n512_));
  AOI21_X1  g390(.A(new_n179_), .B1(new_n178_), .B2(new_n172_), .ZN(new_n513_));
  OAI21_X1  g391(.A(new_n182_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g392(.A1(new_n514_), .A2(G472), .ZN(new_n515_));
  NAND3_X1  g393(.A1(new_n181_), .A2(new_n123_), .A3(new_n182_), .ZN(new_n516_));
  AND4_X1   g394(.A1(KEYINPUT34), .A2(new_n515_), .A3(new_n510_), .A4(new_n516_), .ZN(new_n517_));
  OAI211_X1 g395(.A(new_n389_), .B(new_n324_), .C1(new_n511_), .C2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g396(.A(KEYINPUT35), .B1(new_n470_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n520_));
  INV_X1    g398(.A(new_n518_), .ZN(new_n521_));
  NAND3_X1  g399(.A1(new_n465_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g400(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g401(.A(new_n523_), .B(G110), .ZN(G12));
  AOI22_X1  g402(.A1(new_n515_), .A2(new_n516_), .B1(new_n228_), .B2(new_n509_), .ZN(new_n525_));
  AND2_X1   g403(.A1(new_n389_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g404(.A1(new_n465_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g405(.A1(new_n124_), .A2(G900), .ZN(new_n528_));
  NAND2_X1  g406(.A1(new_n320_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g407(.A1(new_n319_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g408(.A1(new_n501_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g409(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g410(.A(new_n532_), .B(G128), .ZN(G30));
  XNOR2_X1  g411(.A(new_n474_), .B(KEYINPUT36), .ZN(new_n534_));
  NAND2_X1  g412(.A1(new_n175_), .A2(G472), .ZN(new_n535_));
  OR2_X1    g413(.A1(new_n178_), .A2(KEYINPUT37), .ZN(new_n536_));
  NAND3_X1  g414(.A1(new_n178_), .A2(KEYINPUT37), .A3(new_n172_), .ZN(new_n537_));
  NAND2_X1  g415(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g416(.A(new_n535_), .B1(new_n538_), .B2(new_n179_), .ZN(new_n539_));
  NOR2_X1   g417(.A1(new_n123_), .A2(new_n182_), .ZN(new_n540_));
  NOR3_X1   g418(.A1(new_n539_), .A2(new_n184_), .A3(new_n540_), .ZN(new_n541_));
  OAI21_X1  g419(.A(new_n278_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n542_));
  NOR2_X1   g420(.A1(new_n263_), .A2(KEYINPUT25), .ZN(new_n543_));
  OAI21_X1  g421(.A(new_n280_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g422(.A1(new_n284_), .A2(G475), .ZN(new_n545_));
  NAND2_X1  g423(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g424(.A1(new_n546_), .A2(new_n500_), .ZN(new_n547_));
  INV_X1    g425(.A(new_n530_), .ZN(new_n548_));
  NOR2_X1   g426(.A1(new_n326_), .A2(new_n462_), .ZN(new_n549_));
  NAND2_X1  g427(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR4_X1   g428(.A1(new_n541_), .A2(new_n547_), .A3(new_n510_), .A4(new_n550_), .ZN(new_n551_));
  NAND3_X1  g429(.A1(new_n534_), .A2(new_n447_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n553_));
  NAND2_X1  g431(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g432(.A1(new_n534_), .A2(new_n551_), .A3(KEYINPUT38), .A4(new_n447_), .ZN(new_n555_));
  NAND2_X1  g433(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g434(.A(new_n556_), .B(G143), .ZN(G45));
  INV_X1    g435(.A(new_n483_), .ZN(new_n558_));
  NAND2_X1  g436(.A1(new_n558_), .A2(new_n546_), .ZN(new_n559_));
  NOR2_X1   g437(.A1(new_n559_), .A2(new_n530_), .ZN(new_n560_));
  NAND2_X1  g438(.A1(new_n527_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g439(.A(new_n561_), .B(G146), .ZN(G48));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n563_));
  NAND2_X1  g441(.A1(new_n435_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g442(.A(G469), .B1(new_n454_), .B2(G902), .ZN(new_n565_));
  NAND4_X1  g443(.A1(new_n433_), .A2(KEYINPUT39), .A3(new_n434_), .A4(new_n182_), .ZN(new_n566_));
  NAND4_X1  g444(.A1(new_n564_), .A2(new_n448_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g445(.A(new_n236_), .ZN(new_n568_));
  NOR3_X1   g446(.A1(new_n567_), .A2(new_n486_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g447(.A(new_n569_), .B(new_n165_), .ZN(G15));
  INV_X1    g448(.A(new_n567_), .ZN(new_n571_));
  NAND3_X1  g449(.A1(new_n571_), .A2(new_n502_), .A3(new_n236_), .ZN(new_n572_));
  XNOR2_X1  g450(.A(new_n572_), .B(G116), .ZN(G18));
  AND3_X1   g451(.A1(new_n324_), .A2(new_n389_), .A3(new_n525_), .ZN(new_n574_));
  NAND2_X1  g452(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g453(.A(new_n575_), .B(G119), .ZN(G21));
  AOI22_X1  g454(.A1(new_n544_), .A2(new_n545_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n577_));
  INV_X1    g455(.A(new_n235_), .ZN(new_n578_));
  NAND3_X1  g456(.A1(new_n185_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NOR2_X1   g457(.A1(new_n492_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g458(.A1(new_n571_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g459(.A(new_n581_), .B(G122), .ZN(G24));
  NAND2_X1  g460(.A1(new_n474_), .A2(new_n485_), .ZN(new_n583_));
  NAND2_X1  g461(.A1(new_n185_), .A2(new_n510_), .ZN(new_n584_));
  INV_X1    g462(.A(KEYINPUT34), .ZN(new_n585_));
  NAND2_X1  g463(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g464(.A(new_n517_), .ZN(new_n587_));
  AOI21_X1  g465(.A(new_n583_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g466(.A1(new_n588_), .A2(new_n560_), .A3(new_n571_), .ZN(new_n589_));
  XNOR2_X1  g467(.A(new_n589_), .B(G125), .ZN(G27));
  NOR2_X1   g468(.A1(new_n474_), .A2(new_n326_), .ZN(new_n591_));
  NAND2_X1  g469(.A1(new_n560_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g470(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g471(.A1(new_n465_), .A2(new_n236_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g472(.A1(new_n594_), .A2(KEYINPUT40), .ZN(new_n595_));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n596_));
  NAND4_X1  g474(.A1(new_n465_), .A2(new_n596_), .A3(new_n236_), .A4(new_n593_), .ZN(new_n597_));
  NAND2_X1  g475(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g476(.A(KEYINPUT41), .B(G131), .Z(new_n599_));
  XNOR2_X1  g477(.A(new_n598_), .B(new_n599_), .ZN(G33));
  AND2_X1   g478(.A1(new_n591_), .A2(new_n236_), .ZN(new_n601_));
  NAND3_X1  g479(.A1(new_n465_), .A2(new_n531_), .A3(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g480(.A(new_n602_), .B(G134), .ZN(G36));
  NAND2_X1  g481(.A1(new_n499_), .A2(new_n558_), .ZN(new_n604_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n605_));
  NAND2_X1  g483(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g484(.A1(new_n499_), .A2(KEYINPUT42), .A3(new_n558_), .ZN(new_n607_));
  NAND4_X1  g485(.A1(new_n606_), .A2(new_n591_), .A3(new_n525_), .A4(new_n607_), .ZN(new_n608_));
  INV_X1    g486(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g487(.A(new_n434_), .B1(new_n431_), .B2(new_n410_), .ZN(new_n610_));
  AND2_X1   g488(.A1(new_n443_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g489(.A(new_n611_), .B1(G469), .B2(G902), .ZN(new_n612_));
  NAND2_X1  g490(.A1(new_n612_), .A2(new_n435_), .ZN(new_n613_));
  NAND3_X1  g491(.A1(new_n613_), .A2(new_n448_), .A3(new_n548_), .ZN(new_n614_));
  INV_X1    g492(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g493(.A1(new_n609_), .A2(new_n615_), .A3(KEYINPUT43), .ZN(new_n616_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n617_));
  OAI21_X1  g495(.A(new_n617_), .B1(new_n608_), .B2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g496(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g497(.A(KEYINPUT44), .B(G137), .ZN(new_n620_));
  XNOR2_X1  g498(.A(new_n619_), .B(new_n620_), .ZN(G39));
  NAND4_X1  g499(.A1(new_n613_), .A2(new_n185_), .A3(new_n235_), .A4(new_n448_), .ZN(new_n622_));
  NOR2_X1   g500(.A1(new_n622_), .A2(new_n592_), .ZN(new_n623_));
  XOR2_X1   g501(.A(KEYINPUT45), .B(G140), .Z(new_n624_));
  XNOR2_X1  g502(.A(new_n623_), .B(new_n624_), .ZN(G42));
  NOR2_X1   g503(.A1(new_n546_), .A2(new_n483_), .ZN(new_n626_));
  NAND4_X1  g504(.A1(new_n541_), .A2(new_n626_), .A3(new_n578_), .A4(new_n549_), .ZN(new_n627_));
  NOR2_X1   g505(.A1(new_n534_), .A2(new_n627_), .ZN(new_n628_));
  AND4_X1   g506(.A1(new_n564_), .A2(new_n628_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n629_));
  NOR3_X1   g507(.A1(new_n629_), .A2(G952), .A3(G953), .ZN(new_n630_));
  INV_X1    g508(.A(new_n319_), .ZN(new_n631_));
  NAND3_X1  g509(.A1(new_n606_), .A2(new_n631_), .A3(new_n607_), .ZN(new_n632_));
  NOR2_X1   g510(.A1(new_n632_), .A2(new_n472_), .ZN(new_n633_));
  NAND3_X1  g511(.A1(new_n633_), .A2(new_n389_), .A3(new_n571_), .ZN(new_n634_));
  NAND3_X1  g512(.A1(new_n634_), .A2(G952), .A3(new_n186_), .ZN(new_n635_));
  XNOR2_X1  g513(.A(new_n635_), .B(KEYINPUT47), .ZN(new_n636_));
  OR3_X1    g514(.A1(new_n534_), .A2(new_n485_), .A3(new_n472_), .ZN(new_n637_));
  NAND2_X1  g515(.A1(new_n586_), .A2(new_n587_), .ZN(new_n638_));
  OAI21_X1  g516(.A(new_n591_), .B1(new_n638_), .B2(new_n236_), .ZN(new_n639_));
  AOI21_X1  g517(.A(new_n632_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g518(.A1(new_n591_), .A2(new_n578_), .A3(new_n631_), .A4(new_n541_), .ZN(new_n641_));
  NAND2_X1  g519(.A1(new_n285_), .A2(new_n483_), .ZN(new_n642_));
  XNOR2_X1  g520(.A(new_n559_), .B(KEYINPUT46), .ZN(new_n643_));
  AOI21_X1  g521(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g522(.A(new_n571_), .B1(new_n640_), .B2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g523(.A1(new_n564_), .A2(new_n462_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n646_));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n647_));
  NOR2_X1   g525(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n613_), .B2(new_n448_), .ZN(new_n649_));
  AOI21_X1  g527(.A(new_n648_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  AND2_X1   g528(.A1(new_n633_), .A2(new_n591_), .ZN(new_n651_));
  AOI21_X1  g529(.A(new_n629_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  AND3_X1   g530(.A1(new_n636_), .A2(new_n645_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g531(.A(new_n520_), .B1(new_n465_), .B2(new_n521_), .ZN(new_n654_));
  AOI211_X1 g532(.A(KEYINPUT35), .B(new_n518_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n655_));
  NOR2_X1   g533(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g534(.A(new_n560_), .B(new_n591_), .C1(new_n511_), .C2(new_n517_), .ZN(new_n657_));
  INV_X1    g535(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g536(.A1(new_n465_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g537(.A1(new_n389_), .A2(new_n323_), .A3(new_n471_), .A4(new_n577_), .ZN(new_n660_));
  NAND3_X1  g538(.A1(new_n324_), .A2(new_n389_), .A3(new_n525_), .ZN(new_n661_));
  AOI21_X1  g539(.A(new_n567_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g540(.A1(new_n662_), .A2(new_n569_), .ZN(new_n663_));
  NAND4_X1  g541(.A1(new_n659_), .A2(new_n663_), .A3(new_n572_), .A4(new_n589_), .ZN(new_n664_));
  NOR2_X1   g542(.A1(new_n656_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n666_));
  NAND3_X1  g544(.A1(new_n465_), .A2(new_n666_), .A3(new_n548_), .ZN(new_n667_));
  AND2_X1   g545(.A1(new_n591_), .A2(new_n525_), .ZN(new_n668_));
  NOR2_X1   g546(.A1(new_n546_), .A2(new_n500_), .ZN(new_n669_));
  XNOR2_X1  g547(.A(new_n669_), .B(KEYINPUT50), .ZN(new_n670_));
  NOR3_X1   g548(.A1(new_n541_), .A2(new_n547_), .A3(new_n510_), .ZN(new_n671_));
  AOI22_X1  g549(.A1(new_n668_), .A2(new_n670_), .B1(new_n671_), .B2(new_n389_), .ZN(new_n672_));
  OAI21_X1  g550(.A(new_n548_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n673_));
  AOI21_X1  g551(.A(new_n672_), .B1(new_n673_), .B2(KEYINPUT49), .ZN(new_n674_));
  AOI22_X1  g552(.A1(new_n667_), .A2(new_n674_), .B1(new_n452_), .B2(new_n467_), .ZN(new_n675_));
  INV_X1    g553(.A(new_n602_), .ZN(new_n676_));
  AOI21_X1  g554(.A(new_n676_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n677_));
  OAI211_X1 g555(.A(new_n465_), .B(new_n471_), .C1(new_n487_), .C2(new_n502_), .ZN(new_n678_));
  OAI211_X1 g556(.A(new_n465_), .B(new_n526_), .C1(new_n531_), .C2(new_n560_), .ZN(new_n679_));
  AND2_X1   g557(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g558(.A1(new_n665_), .A2(new_n675_), .A3(new_n677_), .A4(new_n680_), .ZN(new_n681_));
  INV_X1    g559(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g560(.A(new_n630_), .B1(new_n653_), .B2(new_n682_), .ZN(G75));
  AND2_X1   g561(.A1(new_n681_), .A2(G902), .ZN(new_n684_));
  INV_X1    g562(.A(new_n377_), .ZN(new_n685_));
  AOI21_X1  g563(.A(new_n371_), .B1(new_n376_), .B2(new_n375_), .ZN(new_n686_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n687_));
  NOR3_X1   g565(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  NAND3_X1  g566(.A1(new_n684_), .A2(new_n328_), .A3(new_n688_), .ZN(new_n689_));
  OR2_X1    g567(.A1(new_n186_), .A2(G952), .ZN(new_n690_));
  NAND2_X1  g568(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g569(.A(new_n688_), .B1(new_n684_), .B2(new_n328_), .ZN(new_n692_));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g571(.A(new_n692_), .ZN(new_n694_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n695_));
  NAND4_X1  g573(.A1(new_n694_), .A2(new_n695_), .A3(new_n690_), .A4(new_n689_), .ZN(new_n696_));
  NAND2_X1  g574(.A1(new_n693_), .A2(new_n696_), .ZN(G51));
  NAND3_X1  g575(.A1(new_n681_), .A2(G469), .A3(G902), .ZN(new_n698_));
  NAND2_X1  g576(.A1(new_n698_), .A2(new_n433_), .ZN(new_n699_));
  NAND3_X1  g577(.A1(new_n681_), .A2(G902), .A3(new_n611_), .ZN(new_n700_));
  NAND2_X1  g578(.A1(new_n700_), .A2(KEYINPUT53), .ZN(new_n701_));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n702_));
  NAND4_X1  g580(.A1(new_n681_), .A2(new_n702_), .A3(G902), .A4(new_n611_), .ZN(new_n703_));
  NAND3_X1  g581(.A1(new_n699_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g582(.A1(new_n704_), .A2(new_n690_), .ZN(new_n705_));
  NAND2_X1  g583(.A1(new_n705_), .A2(KEYINPUT54), .ZN(new_n706_));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n707_));
  NAND3_X1  g585(.A1(new_n704_), .A2(new_n707_), .A3(new_n690_), .ZN(new_n708_));
  NAND2_X1  g586(.A1(new_n706_), .A2(new_n708_), .ZN(G54));
  NOR3_X1   g587(.A1(new_n682_), .A2(new_n493_), .A3(new_n182_), .ZN(new_n710_));
  OR2_X1    g588(.A1(new_n710_), .A2(new_n279_), .ZN(new_n711_));
  NAND2_X1  g589(.A1(new_n710_), .A2(new_n279_), .ZN(new_n712_));
  AND3_X1   g590(.A1(new_n711_), .A2(new_n690_), .A3(new_n712_), .ZN(G60));
  NAND2_X1  g591(.A1(new_n684_), .A2(G478), .ZN(new_n714_));
  INV_X1    g592(.A(new_n481_), .ZN(new_n715_));
  OAI21_X1  g593(.A(new_n690_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g594(.A(new_n716_), .B1(new_n715_), .B2(new_n714_), .ZN(G63));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n718_));
  NAND2_X1  g596(.A1(new_n221_), .A2(new_n224_), .ZN(new_n719_));
  INV_X1    g597(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g598(.A1(new_n684_), .A2(G217), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g599(.A1(new_n721_), .A2(new_n690_), .ZN(new_n722_));
  AOI21_X1  g600(.A(new_n720_), .B1(new_n684_), .B2(G217), .ZN(new_n723_));
  OAI21_X1  g601(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g602(.A(new_n723_), .ZN(new_n725_));
  NAND4_X1  g603(.A1(new_n725_), .A2(KEYINPUT55), .A3(new_n690_), .A4(new_n721_), .ZN(new_n726_));
  NAND2_X1  g604(.A1(new_n724_), .A2(new_n726_), .ZN(G66));
  OAI21_X1  g605(.A(new_n571_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n728_));
  NAND3_X1  g606(.A1(new_n571_), .A2(new_n487_), .A3(new_n236_), .ZN(new_n729_));
  NAND3_X1  g607(.A1(new_n728_), .A2(new_n729_), .A3(new_n572_), .ZN(new_n730_));
  NAND2_X1  g608(.A1(new_n730_), .A2(KEYINPUT56), .ZN(new_n731_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n732_));
  NAND3_X1  g610(.A1(new_n663_), .A2(new_n732_), .A3(new_n572_), .ZN(new_n733_));
  NAND2_X1  g611(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g612(.A1(new_n734_), .A2(new_n468_), .A3(new_n523_), .A4(new_n678_), .ZN(new_n735_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n736_));
  NAND2_X1  g614(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OR2_X1    g615(.A1(new_n492_), .A2(new_n501_), .ZN(new_n738_));
  AOI221_X4 g616(.A(new_n472_), .B1(new_n738_), .B2(new_n486_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n739_));
  AOI21_X1  g617(.A(new_n739_), .B1(new_n522_), .B2(new_n519_), .ZN(new_n740_));
  NAND4_X1  g618(.A1(new_n740_), .A2(KEYINPUT57), .A3(new_n468_), .A4(new_n734_), .ZN(new_n741_));
  NAND3_X1  g619(.A1(new_n737_), .A2(new_n124_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n743_));
  NAND2_X1  g621(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g622(.A1(new_n737_), .A2(KEYINPUT58), .A3(new_n741_), .A4(new_n124_), .ZN(new_n745_));
  NAND2_X1  g623(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g624(.A(new_n356_), .B(new_n370_), .C1(G898), .C2(new_n186_), .ZN(new_n747_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n748_));
  AND2_X1   g626(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g627(.A1(new_n746_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g628(.A(new_n747_), .B(KEYINPUT59), .ZN(new_n751_));
  NAND3_X1  g629(.A1(new_n744_), .A2(new_n745_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g630(.A(new_n124_), .B1(G224), .B2(G898), .ZN(new_n753_));
  INV_X1    g631(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g632(.A1(new_n750_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g633(.A1(new_n747_), .A2(new_n753_), .ZN(new_n756_));
  XNOR2_X1  g634(.A(new_n756_), .B(KEYINPUT60), .ZN(new_n757_));
  NAND2_X1  g635(.A1(new_n755_), .A2(new_n757_), .ZN(G69));
  AOI21_X1  g636(.A(new_n528_), .B1(new_n176_), .B2(new_n199_), .ZN(new_n759_));
  OAI21_X1  g637(.A(new_n759_), .B1(new_n176_), .B2(new_n199_), .ZN(new_n760_));
  INV_X1    g638(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g639(.A(new_n623_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n762_));
  NAND3_X1  g640(.A1(new_n677_), .A2(KEYINPUT61), .A3(new_n762_), .ZN(new_n763_));
  NAND4_X1  g641(.A1(new_n615_), .A2(new_n236_), .A3(new_n389_), .A4(new_n577_), .ZN(new_n764_));
  AND2_X1   g642(.A1(new_n764_), .A2(new_n589_), .ZN(new_n765_));
  NAND3_X1  g643(.A1(new_n763_), .A2(new_n679_), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g644(.A(KEYINPUT61), .B1(new_n677_), .B2(new_n762_), .ZN(new_n767_));
  NOR2_X1   g645(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g646(.A(new_n761_), .B1(new_n768_), .B2(G953), .ZN(new_n769_));
  AND3_X1   g647(.A1(new_n588_), .A2(new_n560_), .A3(new_n571_), .ZN(new_n770_));
  AOI21_X1  g648(.A(new_n770_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n771_));
  AOI21_X1  g649(.A(new_n530_), .B1(new_n643_), .B2(new_n501_), .ZN(new_n772_));
  NAND3_X1  g650(.A1(new_n772_), .A2(new_n465_), .A3(new_n601_), .ZN(new_n773_));
  AND4_X1   g651(.A1(new_n679_), .A2(new_n771_), .A3(new_n762_), .A4(new_n773_), .ZN(new_n774_));
  INV_X1    g652(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g653(.A1(new_n775_), .A2(new_n186_), .A3(new_n760_), .ZN(new_n776_));
  NAND2_X1  g654(.A1(new_n769_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g655(.A(new_n186_), .B1(G227), .B2(G900), .ZN(new_n778_));
  INV_X1    g656(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g657(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g658(.A1(new_n769_), .A2(new_n778_), .A3(new_n776_), .ZN(new_n781_));
  NAND2_X1  g659(.A1(new_n780_), .A2(new_n781_), .ZN(G72));
  INV_X1    g660(.A(new_n730_), .ZN(new_n783_));
  NAND4_X1  g661(.A1(new_n774_), .A2(new_n468_), .A3(new_n783_), .A4(new_n740_), .ZN(new_n784_));
  XNOR2_X1  g662(.A(new_n540_), .B(KEYINPUT62), .ZN(new_n785_));
  AOI21_X1  g663(.A(new_n538_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g664(.A1(new_n681_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n787_));
  AOI21_X1  g665(.A(new_n786_), .B1(KEYINPUT63), .B2(new_n787_), .ZN(new_n788_));
  OR2_X1    g666(.A1(new_n787_), .A2(KEYINPUT63), .ZN(new_n789_));
  AOI21_X1  g667(.A(new_n139_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g668(.A1(new_n538_), .A2(new_n785_), .ZN(new_n791_));
  NAND2_X1  g669(.A1(new_n737_), .A2(new_n741_), .ZN(new_n792_));
  AOI21_X1  g670(.A(new_n791_), .B1(new_n768_), .B2(new_n792_), .ZN(new_n793_));
  AND2_X1   g671(.A1(new_n681_), .A2(new_n540_), .ZN(new_n794_));
  OAI21_X1  g672(.A(new_n139_), .B1(new_n794_), .B2(new_n538_), .ZN(new_n795_));
  OAI21_X1  g673(.A(new_n690_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g674(.A1(new_n790_), .A2(new_n796_), .ZN(G57));
endmodule


