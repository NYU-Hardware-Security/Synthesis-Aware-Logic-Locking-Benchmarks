//Secret key is'0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_c2670" written by ABC on Sun Nov 20 19:50:24 2022

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14,
    G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32,
    G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52,
    G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68,
    G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101,
    G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115,
    G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129,
    G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169,
    G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189,
    G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
    G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213,
    G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248,
    G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264,
    G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276,
    G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860, G868,
    G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981,
    G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096,
    G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446,
    G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445_, new_n447_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n457_, new_n458_, new_n459_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n540_,
    new_n541_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n557_, new_n558_, new_n559_, new_n560_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n586_, new_n587_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1113_, new_n1114_, new_n1115_;
  XOR2_X1   g000(.A(KEYINPUT0), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT1), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  INV_X1    g010(.A(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT3), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT4), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445_));
  XOR2_X1   g020(.A(new_n445_), .B(KEYINPUT5), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447_));
  XNOR2_X1  g022(.A(new_n447_), .B(KEYINPUT6), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n451_));
  XNOR2_X1  g026(.A(new_n451_), .B(KEYINPUT7), .ZN(new_n452_));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453_));
  INV_X1    g028(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g029(.A1(new_n452_), .A2(new_n454_), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452_), .A2(G567), .ZN(new_n457_));
  NAND2_X1  g032(.A1(new_n454_), .A2(G2106), .ZN(new_n458_));
  NAND2_X1  g033(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g034(.A(new_n459_), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461_));
  NAND2_X1  g036(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n462_));
  INV_X1    g037(.A(KEYINPUT9), .ZN(new_n463_));
  NAND2_X1  g038(.A1(new_n463_), .A2(G2104), .ZN(new_n464_));
  NAND2_X1  g039(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g040(.A1(new_n465_), .A2(G125), .A3(G2105), .ZN(new_n466_));
  INV_X1    g041(.A(KEYINPUT10), .ZN(new_n467_));
  NAND2_X1  g042(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g043(.A(G101), .ZN(new_n469_));
  OR2_X1    g044(.A1(KEYINPUT8), .A2(G2105), .ZN(new_n470_));
  NAND2_X1  g045(.A1(KEYINPUT8), .A2(G2105), .ZN(new_n471_));
  AOI21_X1  g046(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g047(.A1(G113), .A2(G2105), .ZN(new_n473_));
  INV_X1    g048(.A(new_n473_), .ZN(new_n474_));
  OAI21_X1  g049(.A(G2104), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g050(.A1(new_n470_), .A2(new_n471_), .ZN(new_n476_));
  NAND3_X1  g051(.A1(new_n476_), .A2(new_n465_), .A3(G137), .ZN(new_n477_));
  INV_X1    g052(.A(G2105), .ZN(new_n478_));
  AOI21_X1  g053(.A(new_n478_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n479_));
  NAND3_X1  g054(.A1(new_n479_), .A2(KEYINPUT10), .A3(G125), .ZN(new_n480_));
  NAND4_X1  g055(.A1(new_n468_), .A2(new_n475_), .A3(new_n477_), .A4(new_n480_), .ZN(new_n481_));
  INV_X1    g056(.A(new_n481_), .ZN(G160));
  AND2_X1   g057(.A1(KEYINPUT8), .A2(G2105), .ZN(new_n483_));
  NOR2_X1   g058(.A1(KEYINPUT8), .A2(G2105), .ZN(new_n484_));
  NOR2_X1   g059(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g060(.A1(new_n485_), .A2(new_n461_), .ZN(new_n486_));
  AOI22_X1  g061(.A1(new_n462_), .A2(new_n464_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n487_));
  AOI22_X1  g062(.A1(G100), .A2(new_n486_), .B1(new_n487_), .B2(G136), .ZN(new_n488_));
  AOI22_X1  g063(.A1(new_n465_), .A2(G124), .B1(G112), .B2(G2104), .ZN(new_n489_));
  OAI21_X1  g064(.A(new_n488_), .B1(new_n478_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g065(.A(new_n490_), .B(KEYINPUT11), .ZN(new_n491_));
  XNOR2_X1  g066(.A(new_n491_), .B(KEYINPUT12), .ZN(G162));
  XNOR2_X1  g067(.A(KEYINPUT9), .B(G2104), .ZN(new_n493_));
  OAI21_X1  g068(.A(G138), .B1(new_n483_), .B2(new_n484_), .ZN(new_n494_));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495_));
  AOI21_X1  g070(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g071(.A(G102), .B1(new_n483_), .B2(new_n484_), .ZN(new_n497_));
  NAND2_X1  g072(.A1(G114), .A2(G2105), .ZN(new_n498_));
  AOI21_X1  g073(.A(new_n461_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g074(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g075(.A(new_n500_), .B(KEYINPUT13), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502_));
  NAND3_X1  g077(.A1(new_n502_), .A2(G50), .A3(G543), .ZN(new_n503_));
  XOR2_X1   g078(.A(new_n503_), .B(KEYINPUT14), .Z(new_n504_));
  NOR2_X1   g079(.A1(G543), .A2(G651), .ZN(new_n505_));
  NAND2_X1  g080(.A1(new_n505_), .A2(G88), .ZN(new_n506_));
  INV_X1    g081(.A(G543), .ZN(new_n507_));
  NOR2_X1   g082(.A1(new_n507_), .A2(G75), .ZN(new_n508_));
  OAI21_X1  g083(.A(G651), .B1(G62), .B2(G543), .ZN(new_n509_));
  OAI211_X1 g084(.A(new_n504_), .B(new_n506_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g085(.A(KEYINPUT15), .ZN(new_n511_));
  OR2_X1    g086(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g087(.A1(new_n510_), .A2(new_n511_), .ZN(new_n513_));
  NAND2_X1  g088(.A1(new_n512_), .A2(new_n513_), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(new_n502_), .A2(G51), .A3(G543), .ZN(new_n516_));
  XOR2_X1   g091(.A(new_n516_), .B(KEYINPUT17), .Z(new_n517_));
  NOR2_X1   g092(.A1(new_n507_), .A2(G76), .ZN(new_n518_));
  OAI21_X1  g093(.A(G651), .B1(G63), .B2(G543), .ZN(new_n519_));
  OAI21_X1  g094(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g095(.A1(new_n505_), .A2(G89), .ZN(new_n521_));
  XOR2_X1   g096(.A(new_n521_), .B(KEYINPUT16), .Z(new_n522_));
  OR2_X1    g097(.A1(new_n520_), .A2(new_n522_), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  OR2_X1    g099(.A1(G64), .A2(G543), .ZN(new_n525_));
  OAI211_X1 g100(.A(new_n525_), .B(G651), .C1(G77), .C2(new_n507_), .ZN(new_n526_));
  OR2_X1    g101(.A1(G90), .A2(G543), .ZN(new_n527_));
  OAI211_X1 g102(.A(new_n527_), .B(new_n502_), .C1(G52), .C2(new_n507_), .ZN(new_n528_));
  NAND2_X1  g103(.A1(new_n526_), .A2(new_n528_), .ZN(G301));
  INV_X1    g104(.A(G301), .ZN(G171));
  AOI21_X1  g105(.A(new_n502_), .B1(G56), .B2(new_n507_), .ZN(new_n531_));
  INV_X1    g106(.A(G68), .ZN(new_n532_));
  OAI21_X1  g107(.A(new_n531_), .B1(new_n532_), .B2(new_n507_), .ZN(new_n533_));
  AOI21_X1  g108(.A(G651), .B1(new_n507_), .B2(G81), .ZN(new_n534_));
  INV_X1    g109(.A(G43), .ZN(new_n535_));
  OAI21_X1  g110(.A(new_n534_), .B1(new_n535_), .B2(new_n507_), .ZN(new_n536_));
  NAND2_X1  g111(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g112(.A1(new_n537_), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540_));
  NAND4_X1  g115(.A1(G319), .A2(G483), .A3(G661), .A4(new_n540_), .ZN(new_n541_));
  XOR2_X1   g116(.A(new_n541_), .B(KEYINPUT18), .Z(G188));
  OAI21_X1  g117(.A(G651), .B1(G65), .B2(G543), .ZN(new_n543_));
  INV_X1    g118(.A(G78), .ZN(new_n544_));
  AOI21_X1  g119(.A(new_n543_), .B1(new_n544_), .B2(G543), .ZN(new_n545_));
  OR2_X1    g120(.A1(new_n507_), .A2(G53), .ZN(new_n546_));
  INV_X1    g121(.A(G91), .ZN(new_n547_));
  AOI21_X1  g122(.A(G651), .B1(new_n547_), .B2(new_n507_), .ZN(new_n548_));
  AOI21_X1  g123(.A(new_n545_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g124(.A(new_n549_), .ZN(G299));
  AOI21_X1  g125(.A(G651), .B1(new_n507_), .B2(G87), .ZN(new_n551_));
  INV_X1    g126(.A(G49), .ZN(new_n552_));
  OAI21_X1  g127(.A(new_n551_), .B1(new_n552_), .B2(new_n507_), .ZN(new_n553_));
  OR2_X1    g128(.A1(new_n507_), .A2(G74), .ZN(new_n554_));
  OAI21_X1  g129(.A(new_n553_), .B1(new_n502_), .B2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g130(.A(new_n555_), .B(KEYINPUT19), .Z(G288));
  OR2_X1    g131(.A1(G61), .A2(G543), .ZN(new_n557_));
  OAI211_X1 g132(.A(new_n557_), .B(G651), .C1(G73), .C2(new_n507_), .ZN(new_n558_));
  OR2_X1    g133(.A1(G86), .A2(G543), .ZN(new_n559_));
  OAI211_X1 g134(.A(new_n559_), .B(new_n502_), .C1(G48), .C2(new_n507_), .ZN(new_n560_));
  NAND2_X1  g135(.A1(new_n558_), .A2(new_n560_), .ZN(G305));
  NAND3_X1  g136(.A1(new_n502_), .A2(G47), .A3(G543), .ZN(new_n562_));
  XOR2_X1   g137(.A(new_n562_), .B(KEYINPUT21), .Z(new_n563_));
  NAND2_X1  g138(.A1(new_n505_), .A2(G85), .ZN(new_n564_));
  XNOR2_X1  g139(.A(new_n564_), .B(KEYINPUT20), .ZN(new_n565_));
  NAND3_X1  g140(.A1(G72), .A2(G543), .A3(G651), .ZN(new_n566_));
  NAND3_X1  g141(.A1(new_n507_), .A2(G60), .A3(G651), .ZN(new_n567_));
  XNOR2_X1  g142(.A(new_n567_), .B(KEYINPUT22), .ZN(new_n568_));
  NAND4_X1  g143(.A1(new_n563_), .A2(new_n565_), .A3(new_n566_), .A4(new_n568_), .ZN(G290));
  NAND2_X1  g144(.A1(G301), .A2(G868), .ZN(new_n570_));
  NAND3_X1  g145(.A1(new_n502_), .A2(G54), .A3(G543), .ZN(new_n571_));
  INV_X1    g146(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g147(.A1(G66), .A2(G543), .ZN(new_n573_));
  OAI211_X1 g148(.A(new_n573_), .B(G651), .C1(G79), .C2(new_n507_), .ZN(new_n574_));
  INV_X1    g149(.A(G92), .ZN(new_n575_));
  INV_X1    g150(.A(new_n505_), .ZN(new_n576_));
  OAI21_X1  g151(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n578_));
  NAND2_X1  g153(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g154(.A(new_n574_), .B(KEYINPUT23), .C1(new_n575_), .C2(new_n576_), .ZN(new_n580_));
  AOI21_X1  g155(.A(new_n572_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g156(.A(new_n581_), .B(KEYINPUT24), .ZN(new_n582_));
  INV_X1    g157(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g158(.A(new_n570_), .B1(new_n583_), .B2(G868), .ZN(G284));
  XNOR2_X1  g159(.A(G284), .B(KEYINPUT25), .ZN(G321));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G868), .ZN(new_n586_));
  NAND2_X1  g161(.A1(G299), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g162(.A(new_n587_), .B1(G168), .B2(new_n586_), .ZN(G297));
  OAI21_X1  g163(.A(new_n587_), .B1(G168), .B2(new_n586_), .ZN(G280));
  INV_X1    g164(.A(G559), .ZN(new_n590_));
  AOI21_X1  g165(.A(G860), .B1(new_n590_), .B2(KEYINPUT27), .ZN(new_n591_));
  OAI21_X1  g166(.A(new_n591_), .B1(KEYINPUT27), .B2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g167(.A1(new_n583_), .A2(new_n592_), .ZN(G148));
  INV_X1    g168(.A(new_n537_), .ZN(new_n594_));
  NAND2_X1  g169(.A1(new_n594_), .A2(new_n586_), .ZN(new_n595_));
  INV_X1    g170(.A(new_n581_), .ZN(new_n596_));
  NOR2_X1   g171(.A1(new_n596_), .A2(G559), .ZN(new_n597_));
  OAI21_X1  g172(.A(new_n595_), .B1(new_n597_), .B2(new_n586_), .ZN(G282));
  OAI21_X1  g173(.A(new_n595_), .B1(new_n597_), .B2(new_n586_), .ZN(G323));
  AOI22_X1  g174(.A1(G99), .A2(new_n486_), .B1(new_n487_), .B2(G135), .ZN(new_n600_));
  NAND3_X1  g175(.A1(G111), .A2(G2104), .A3(G2105), .ZN(new_n601_));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n602_));
  OR2_X1    g177(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g178(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  AOI22_X1  g179(.A1(G123), .A2(new_n479_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g180(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g181(.A(new_n606_), .B(KEYINPUT29), .Z(new_n607_));
  XOR2_X1   g182(.A(new_n607_), .B(G2096), .Z(new_n608_));
  OAI21_X1  g183(.A(new_n486_), .B1(new_n463_), .B2(G2105), .ZN(new_n609_));
  XOR2_X1   g184(.A(new_n609_), .B(G2100), .Z(new_n610_));
  NAND2_X1  g185(.A1(new_n608_), .A2(new_n610_), .ZN(G156));
  XNOR2_X1  g186(.A(G2427), .B(G2430), .ZN(new_n612_));
  XNOR2_X1  g187(.A(G2435), .B(G2438), .ZN(new_n613_));
  OR2_X1    g188(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g189(.A(G2443), .B(G2446), .ZN(new_n615_));
  NOR2_X1   g190(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g191(.A(new_n616_), .B(KEYINPUT30), .ZN(new_n617_));
  NAND2_X1  g192(.A1(new_n612_), .A2(new_n613_), .ZN(new_n618_));
  NOR2_X1   g193(.A1(new_n618_), .A2(new_n615_), .ZN(new_n619_));
  XNOR2_X1  g194(.A(new_n619_), .B(KEYINPUT31), .ZN(new_n620_));
  NAND3_X1  g195(.A1(new_n614_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n621_));
  NAND3_X1  g196(.A1(new_n617_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g197(.A(KEYINPUT32), .B(G2451), .ZN(new_n623_));
  XOR2_X1   g198(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625_));
  XNOR2_X1  g200(.A(KEYINPUT33), .B(G2454), .ZN(new_n626_));
  XOR2_X1   g201(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  INV_X1    g202(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g203(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g204(.A(new_n622_), .B(new_n623_), .ZN(new_n630_));
  NAND2_X1  g205(.A1(new_n630_), .A2(new_n627_), .ZN(new_n631_));
  NAND3_X1  g206(.A1(new_n629_), .A2(G14), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g207(.A(new_n632_), .ZN(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634_));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635_));
  INV_X1    g210(.A(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637_));
  OR2_X1    g212(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g213(.A(KEYINPUT35), .ZN(new_n639_));
  AOI21_X1  g214(.A(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g215(.A(new_n638_), .ZN(new_n641_));
  NOR2_X1   g216(.A1(new_n641_), .A2(KEYINPUT34), .ZN(new_n642_));
  NAND2_X1  g217(.A1(new_n636_), .A2(new_n637_), .ZN(new_n643_));
  AOI21_X1  g218(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  MUX2_X1   g219(.A(new_n640_), .B(new_n634_), .S(new_n644_), .Z(new_n645_));
  XNOR2_X1  g220(.A(KEYINPUT36), .B(KEYINPUT37), .ZN(new_n646_));
  XNOR2_X1  g221(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g222(.A(G2096), .B(G2100), .ZN(new_n648_));
  XOR2_X1   g223(.A(new_n647_), .B(new_n648_), .Z(G227));
  XNOR2_X1  g224(.A(G1961), .B(G1966), .ZN(new_n650_));
  INV_X1    g225(.A(KEYINPUT38), .ZN(new_n651_));
  XNOR2_X1  g226(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g227(.A(G1956), .B(G2474), .ZN(new_n653_));
  NAND2_X1  g228(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655_));
  XNOR2_X1  g230(.A(new_n655_), .B(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g231(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g232(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g233(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND2_X1  g234(.A1(new_n654_), .A2(new_n656_), .ZN(new_n660_));
  NOR2_X1   g235(.A1(new_n652_), .A2(new_n653_), .ZN(new_n661_));
  MUX2_X1   g236(.A(new_n660_), .B(new_n656_), .S(new_n661_), .Z(new_n662_));
  NAND2_X1  g237(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664_));
  XNOR2_X1  g239(.A(KEYINPUT41), .B(KEYINPUT42), .ZN(new_n665_));
  XNOR2_X1  g240(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g241(.A(new_n663_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668_));
  OR2_X1    g243(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g244(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NAND2_X1  g245(.A1(new_n669_), .A2(new_n670_), .ZN(G229));
  MUX2_X1   g246(.A(G35), .B(new_n491_), .S(G29), .Z(new_n672_));
  XNOR2_X1  g247(.A(KEYINPUT66), .B(G2090), .ZN(new_n673_));
  XOR2_X1   g248(.A(new_n672_), .B(new_n673_), .Z(new_n674_));
  INV_X1    g249(.A(new_n674_), .ZN(new_n675_));
  AND2_X1   g250(.A1(new_n675_), .A2(KEYINPUT67), .ZN(new_n676_));
  NOR2_X1   g251(.A1(new_n675_), .A2(KEYINPUT67), .ZN(new_n677_));
  INV_X1    g252(.A(G29), .ZN(new_n678_));
  AND2_X1   g253(.A1(new_n678_), .A2(G33), .ZN(new_n679_));
  NAND2_X1  g254(.A1(new_n486_), .A2(G103), .ZN(new_n680_));
  NAND2_X1  g255(.A1(new_n487_), .A2(G139), .ZN(new_n681_));
  NAND2_X1  g256(.A1(new_n479_), .A2(G127), .ZN(new_n682_));
  NAND3_X1  g257(.A1(G115), .A2(G2104), .A3(G2105), .ZN(new_n683_));
  XNOR2_X1  g258(.A(new_n683_), .B(KEYINPUT56), .ZN(new_n684_));
  NAND4_X1  g259(.A1(new_n680_), .A2(new_n681_), .A3(new_n682_), .A4(new_n684_), .ZN(new_n685_));
  AOI21_X1  g260(.A(new_n679_), .B1(new_n685_), .B2(G29), .ZN(new_n686_));
  XOR2_X1   g261(.A(KEYINPUT57), .B(G2072), .Z(new_n687_));
  NOR2_X1   g262(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g263(.A(G16), .ZN(new_n689_));
  OAI21_X1  g264(.A(new_n689_), .B1(KEYINPUT72), .B2(G23), .ZN(new_n690_));
  AOI21_X1  g265(.A(new_n690_), .B1(KEYINPUT72), .B2(G23), .ZN(new_n691_));
  INV_X1    g266(.A(G288), .ZN(new_n692_));
  AOI21_X1  g267(.A(new_n691_), .B1(new_n692_), .B2(G16), .ZN(new_n693_));
  MUX2_X1   g268(.A(G24), .B(G290), .S(G16), .Z(new_n694_));
  OAI22_X1  g269(.A1(new_n693_), .A2(G1976), .B1(G1986), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g270(.A(new_n688_), .B(new_n695_), .C1(G1986), .C2(new_n694_), .ZN(new_n696_));
  AND2_X1   g271(.A1(new_n686_), .A2(new_n687_), .ZN(new_n697_));
  INV_X1    g272(.A(G11), .ZN(new_n698_));
  INV_X1    g273(.A(G868), .ZN(new_n699_));
  AOI21_X1  g274(.A(new_n698_), .B1(KEYINPUT26), .B2(new_n699_), .ZN(new_n700_));
  AND2_X1   g275(.A1(KEYINPUT69), .A2(G28), .ZN(new_n701_));
  OAI21_X1  g276(.A(new_n678_), .B1(KEYINPUT69), .B2(G28), .ZN(new_n702_));
  AND2_X1   g277(.A1(new_n689_), .A2(G6), .ZN(new_n703_));
  AOI21_X1  g278(.A(new_n703_), .B1(G305), .B2(G16), .ZN(new_n704_));
  XNOR2_X1  g279(.A(KEYINPUT70), .B(G1981), .ZN(new_n705_));
  OAI221_X1 g280(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g281(.A(new_n706_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n707_));
  OAI21_X1  g282(.A(new_n707_), .B1(new_n607_), .B2(new_n678_), .ZN(new_n708_));
  AOI211_X1 g283(.A(new_n697_), .B(new_n708_), .C1(G1976), .C2(new_n693_), .ZN(new_n709_));
  INV_X1    g284(.A(G26), .ZN(new_n710_));
  OR3_X1    g285(.A1(new_n710_), .A2(KEYINPUT62), .A3(G29), .ZN(new_n711_));
  OAI21_X1  g286(.A(KEYINPUT62), .B1(new_n710_), .B2(G29), .ZN(new_n712_));
  NAND2_X1  g287(.A1(new_n486_), .A2(G104), .ZN(new_n713_));
  XOR2_X1   g288(.A(new_n713_), .B(KEYINPUT64), .Z(new_n714_));
  NAND2_X1  g289(.A1(new_n476_), .A2(new_n465_), .ZN(new_n715_));
  INV_X1    g290(.A(G140), .ZN(new_n716_));
  OR3_X1    g291(.A1(new_n715_), .A2(KEYINPUT63), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g292(.A(KEYINPUT63), .B1(new_n715_), .B2(new_n716_), .ZN(new_n718_));
  NAND2_X1  g293(.A1(G116), .A2(G2104), .ZN(new_n719_));
  INV_X1    g294(.A(G128), .ZN(new_n720_));
  OAI21_X1  g295(.A(new_n719_), .B1(new_n493_), .B2(new_n720_), .ZN(new_n721_));
  AOI22_X1  g296(.A1(new_n717_), .A2(new_n718_), .B1(G2105), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g297(.A1(new_n714_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g298(.A(new_n723_), .ZN(new_n724_));
  OAI211_X1 g299(.A(new_n711_), .B(new_n712_), .C1(new_n724_), .C2(new_n678_), .ZN(new_n725_));
  XNOR2_X1  g300(.A(KEYINPUT65), .B(G2067), .ZN(new_n726_));
  XNOR2_X1  g301(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g302(.A1(new_n696_), .A2(new_n709_), .A3(new_n727_), .ZN(new_n728_));
  NOR3_X1   g303(.A1(new_n676_), .A2(new_n677_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g304(.A1(new_n689_), .A2(G22), .ZN(new_n730_));
  OAI21_X1  g305(.A(new_n730_), .B1(G166), .B2(new_n689_), .ZN(new_n731_));
  XNOR2_X1  g306(.A(new_n731_), .B(KEYINPUT71), .ZN(new_n732_));
  INV_X1    g307(.A(G1971), .ZN(new_n733_));
  XNOR2_X1  g308(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  NAND2_X1  g309(.A1(new_n678_), .A2(G25), .ZN(new_n735_));
  AOI22_X1  g310(.A1(G95), .A2(new_n486_), .B1(new_n487_), .B2(G131), .ZN(new_n736_));
  AOI22_X1  g311(.A1(new_n465_), .A2(G119), .B1(G107), .B2(G2104), .ZN(new_n737_));
  OAI21_X1  g312(.A(new_n736_), .B1(new_n478_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g313(.A(new_n738_), .B(KEYINPUT73), .ZN(new_n739_));
  INV_X1    g314(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g315(.A(new_n735_), .B1(new_n740_), .B2(new_n678_), .ZN(new_n741_));
  XNOR2_X1  g316(.A(new_n741_), .B(G1991), .ZN(new_n742_));
  NOR2_X1   g317(.A1(G27), .A2(G29), .ZN(new_n743_));
  AOI21_X1  g318(.A(new_n743_), .B1(new_n500_), .B2(G29), .ZN(new_n744_));
  XOR2_X1   g319(.A(KEYINPUT68), .B(G2078), .Z(new_n745_));
  XNOR2_X1  g320(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  AND2_X1   g321(.A1(KEYINPUT58), .A2(G32), .ZN(new_n747_));
  NOR2_X1   g322(.A1(KEYINPUT58), .A2(G32), .ZN(new_n748_));
  OAI21_X1  g323(.A(new_n678_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g324(.A(new_n749_), .B(KEYINPUT59), .ZN(new_n750_));
  NAND2_X1  g325(.A1(new_n487_), .A2(G141), .ZN(new_n751_));
  XNOR2_X1  g326(.A(new_n751_), .B(KEYINPUT60), .ZN(new_n752_));
  NAND2_X1  g327(.A1(G117), .A2(G2104), .ZN(new_n753_));
  INV_X1    g328(.A(G129), .ZN(new_n754_));
  OAI21_X1  g329(.A(new_n753_), .B1(new_n493_), .B2(new_n754_), .ZN(new_n755_));
  AOI22_X1  g330(.A1(new_n755_), .A2(G2105), .B1(new_n486_), .B2(G105), .ZN(new_n756_));
  NAND2_X1  g331(.A1(new_n752_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g332(.A(new_n750_), .B1(new_n757_), .B2(G29), .ZN(new_n758_));
  XOR2_X1   g333(.A(KEYINPUT61), .B(G1996), .Z(new_n759_));
  XNOR2_X1  g334(.A(new_n758_), .B(new_n759_), .ZN(new_n760_));
  NOR4_X1   g335(.A1(new_n734_), .A2(new_n742_), .A3(new_n746_), .A4(new_n760_), .ZN(new_n761_));
  NAND2_X1  g336(.A1(new_n689_), .A2(G5), .ZN(new_n762_));
  OAI21_X1  g337(.A(new_n762_), .B1(G171), .B2(new_n689_), .ZN(new_n763_));
  XOR2_X1   g338(.A(new_n763_), .B(G1961), .Z(new_n764_));
  NAND2_X1  g339(.A1(new_n689_), .A2(G20), .ZN(new_n765_));
  XNOR2_X1  g340(.A(new_n765_), .B(KEYINPUT48), .ZN(new_n766_));
  AOI21_X1  g341(.A(new_n766_), .B1(G299), .B2(G16), .ZN(new_n767_));
  XNOR2_X1  g342(.A(new_n767_), .B(G1956), .ZN(new_n768_));
  NAND2_X1  g343(.A1(new_n689_), .A2(G19), .ZN(new_n769_));
  XOR2_X1   g344(.A(new_n769_), .B(KEYINPUT43), .Z(new_n770_));
  OAI21_X1  g345(.A(new_n770_), .B1(new_n537_), .B2(new_n689_), .ZN(new_n771_));
  XNOR2_X1  g346(.A(new_n771_), .B(KEYINPUT45), .ZN(new_n772_));
  XNOR2_X1  g347(.A(KEYINPUT44), .B(G1341), .ZN(new_n773_));
  INV_X1    g348(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g349(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g350(.A1(new_n764_), .A2(new_n768_), .A3(new_n775_), .ZN(new_n776_));
  XOR2_X1   g351(.A(KEYINPUT47), .B(G1348), .Z(new_n777_));
  INV_X1    g352(.A(new_n777_), .ZN(new_n778_));
  INV_X1    g353(.A(KEYINPUT46), .ZN(new_n779_));
  INV_X1    g354(.A(G4), .ZN(new_n780_));
  AOI21_X1  g355(.A(G16), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g356(.A(new_n781_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n782_));
  OAI21_X1  g357(.A(new_n782_), .B1(new_n596_), .B2(new_n689_), .ZN(new_n783_));
  AOI21_X1  g358(.A(new_n776_), .B1(new_n778_), .B2(new_n783_), .ZN(new_n784_));
  OR2_X1    g359(.A1(new_n772_), .A2(new_n774_), .ZN(new_n785_));
  OR2_X1    g360(.A1(KEYINPUT49), .A2(G21), .ZN(new_n786_));
  NAND2_X1  g361(.A1(KEYINPUT49), .A2(G21), .ZN(new_n787_));
  AOI21_X1  g362(.A(G16), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g363(.A(new_n788_), .B1(G286), .B2(G16), .ZN(new_n789_));
  XNOR2_X1  g364(.A(KEYINPUT50), .B(G1966), .ZN(new_n790_));
  XNOR2_X1  g365(.A(new_n789_), .B(new_n790_), .ZN(new_n791_));
  OR2_X1    g366(.A1(new_n783_), .A2(new_n778_), .ZN(new_n792_));
  NAND4_X1  g367(.A1(new_n784_), .A2(new_n785_), .A3(new_n791_), .A4(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g368(.A(new_n793_), .B(KEYINPUT51), .ZN(new_n794_));
  INV_X1    g369(.A(KEYINPUT52), .ZN(new_n795_));
  OR2_X1    g370(.A1(new_n795_), .A2(G34), .ZN(new_n796_));
  NAND2_X1  g371(.A1(new_n795_), .A2(G34), .ZN(new_n797_));
  AOI21_X1  g372(.A(G29), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g373(.A(new_n798_), .B(KEYINPUT53), .ZN(new_n799_));
  NAND2_X1  g374(.A1(new_n481_), .A2(KEYINPUT54), .ZN(new_n800_));
  OAI21_X1  g375(.A(new_n473_), .B1(new_n485_), .B2(new_n469_), .ZN(new_n801_));
  AOI22_X1  g376(.A1(new_n801_), .A2(G2104), .B1(new_n487_), .B2(G137), .ZN(new_n802_));
  INV_X1    g377(.A(KEYINPUT54), .ZN(new_n803_));
  NAND4_X1  g378(.A1(new_n802_), .A2(new_n803_), .A3(new_n468_), .A4(new_n480_), .ZN(new_n804_));
  AND2_X1   g379(.A1(new_n800_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g380(.A(new_n799_), .B1(new_n805_), .B2(new_n678_), .ZN(new_n806_));
  XNOR2_X1  g381(.A(new_n806_), .B(KEYINPUT55), .ZN(new_n807_));
  INV_X1    g382(.A(G2084), .ZN(new_n808_));
  XNOR2_X1  g383(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  NAND4_X1  g384(.A1(new_n729_), .A2(new_n761_), .A3(new_n794_), .A4(new_n809_), .ZN(G150));
  XNOR2_X1  g385(.A(G150), .B(KEYINPUT74), .ZN(G311));
  NOR2_X1   g386(.A1(KEYINPUT76), .A2(G860), .ZN(new_n812_));
  XNOR2_X1  g387(.A(new_n537_), .B(KEYINPUT77), .ZN(new_n813_));
  NAND3_X1  g388(.A1(new_n813_), .A2(new_n581_), .A3(G559), .ZN(new_n814_));
  INV_X1    g389(.A(G860), .ZN(new_n815_));
  NAND2_X1  g390(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g391(.A(new_n813_), .B1(new_n581_), .B2(G559), .ZN(new_n817_));
  OAI21_X1  g392(.A(KEYINPUT76), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g393(.A1(G80), .A2(G543), .A3(G651), .ZN(new_n819_));
  XOR2_X1   g394(.A(new_n819_), .B(KEYINPUT75), .Z(new_n820_));
  INV_X1    g395(.A(G67), .ZN(new_n821_));
  OAI21_X1  g396(.A(G651), .B1(new_n821_), .B2(G543), .ZN(new_n822_));
  OAI221_X1 g397(.A(new_n822_), .B1(G55), .B2(new_n507_), .C1(new_n576_), .C2(G93), .ZN(new_n823_));
  NAND2_X1  g398(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g399(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g400(.A(new_n812_), .B1(new_n818_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g401(.A(new_n826_), .B1(new_n818_), .B2(new_n825_), .ZN(G145));
  AND2_X1   g402(.A1(new_n752_), .A2(new_n756_), .ZN(new_n828_));
  INV_X1    g403(.A(new_n496_), .ZN(new_n829_));
  NAND2_X1  g404(.A1(new_n497_), .A2(new_n498_), .ZN(new_n830_));
  NAND2_X1  g405(.A1(new_n830_), .A2(G2104), .ZN(new_n831_));
  NAND2_X1  g406(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g407(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g408(.A1(new_n757_), .A2(new_n500_), .ZN(new_n834_));
  NAND3_X1  g409(.A1(new_n833_), .A2(new_n739_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g410(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g411(.A(new_n739_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n837_));
  NOR3_X1   g412(.A1(new_n836_), .A2(new_n837_), .A3(G160), .ZN(new_n838_));
  INV_X1    g413(.A(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g414(.A(new_n723_), .B(KEYINPUT81), .ZN(new_n840_));
  NAND2_X1  g415(.A1(new_n487_), .A2(G142), .ZN(new_n841_));
  XNOR2_X1  g416(.A(new_n841_), .B(KEYINPUT78), .ZN(new_n842_));
  NAND2_X1  g417(.A1(new_n486_), .A2(G106), .ZN(new_n843_));
  INV_X1    g418(.A(KEYINPUT79), .ZN(new_n844_));
  NAND2_X1  g419(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g420(.A1(new_n486_), .A2(KEYINPUT79), .A3(G106), .ZN(new_n846_));
  NAND2_X1  g421(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g422(.A1(G118), .A2(G2104), .A3(G2105), .ZN(new_n848_));
  NAND2_X1  g423(.A1(new_n479_), .A2(G130), .ZN(new_n849_));
  XNOR2_X1  g424(.A(new_n849_), .B(KEYINPUT80), .ZN(new_n850_));
  NAND4_X1  g425(.A1(new_n842_), .A2(new_n847_), .A3(new_n848_), .A4(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g426(.A(new_n851_), .B(new_n685_), .ZN(new_n852_));
  NAND2_X1  g427(.A1(new_n840_), .A2(new_n852_), .ZN(new_n853_));
  OR2_X1    g428(.A1(new_n840_), .A2(new_n852_), .ZN(new_n854_));
  OAI21_X1  g429(.A(G160), .B1(new_n836_), .B2(new_n837_), .ZN(new_n855_));
  NAND4_X1  g430(.A1(new_n839_), .A2(new_n853_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g431(.A1(new_n854_), .A2(new_n853_), .ZN(new_n857_));
  INV_X1    g432(.A(new_n837_), .ZN(new_n858_));
  AOI21_X1  g433(.A(new_n481_), .B1(new_n858_), .B2(new_n835_), .ZN(new_n859_));
  OAI21_X1  g434(.A(new_n857_), .B1(new_n838_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g435(.A1(new_n856_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g436(.A(new_n607_), .B(new_n609_), .ZN(new_n862_));
  XNOR2_X1  g437(.A(new_n491_), .B(KEYINPUT82), .ZN(new_n863_));
  XNOR2_X1  g438(.A(new_n862_), .B(new_n863_), .ZN(new_n864_));
  NAND2_X1  g439(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g440(.A(G37), .ZN(new_n866_));
  INV_X1    g441(.A(new_n864_), .ZN(new_n867_));
  NAND3_X1  g442(.A1(new_n867_), .A2(new_n856_), .A3(new_n860_), .ZN(new_n868_));
  NAND3_X1  g443(.A1(new_n865_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g444(.A(new_n869_), .ZN(G395));
  XNOR2_X1  g445(.A(G288), .B(KEYINPUT87), .ZN(new_n871_));
  XNOR2_X1  g446(.A(G305), .B(KEYINPUT86), .ZN(new_n872_));
  XNOR2_X1  g447(.A(new_n871_), .B(new_n872_), .ZN(new_n873_));
  XOR2_X1   g448(.A(G303), .B(G290), .Z(new_n874_));
  XNOR2_X1  g449(.A(new_n873_), .B(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g450(.A(new_n875_), .B(KEYINPUT85), .ZN(new_n876_));
  XNOR2_X1  g451(.A(new_n581_), .B(G299), .ZN(new_n877_));
  XNOR2_X1  g452(.A(new_n824_), .B(new_n594_), .ZN(new_n878_));
  NAND3_X1  g453(.A1(new_n877_), .A2(new_n597_), .A3(new_n878_), .ZN(new_n879_));
  XOR2_X1   g454(.A(new_n879_), .B(KEYINPUT84), .Z(new_n880_));
  INV_X1    g455(.A(KEYINPUT83), .ZN(new_n881_));
  XNOR2_X1  g456(.A(new_n878_), .B(new_n881_), .ZN(new_n882_));
  INV_X1    g457(.A(new_n877_), .ZN(new_n883_));
  NAND3_X1  g458(.A1(new_n882_), .A2(new_n597_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g459(.A1(new_n882_), .A2(new_n877_), .ZN(new_n885_));
  NAND2_X1  g460(.A1(new_n883_), .A2(new_n878_), .ZN(new_n886_));
  NAND2_X1  g461(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g462(.A(new_n887_), .ZN(new_n888_));
  OAI211_X1 g463(.A(new_n880_), .B(new_n884_), .C1(new_n597_), .C2(new_n888_), .ZN(new_n889_));
  XOR2_X1   g464(.A(new_n876_), .B(new_n889_), .Z(new_n890_));
  MUX2_X1   g465(.A(new_n890_), .B(new_n824_), .S(new_n586_), .Z(G295));
  MUX2_X1   g466(.A(new_n890_), .B(new_n824_), .S(new_n586_), .Z(G331));
  XOR2_X1   g467(.A(new_n873_), .B(new_n874_), .Z(new_n893_));
  NAND2_X1  g468(.A1(new_n882_), .A2(new_n883_), .ZN(new_n894_));
  NAND2_X1  g469(.A1(new_n877_), .A2(new_n878_), .ZN(new_n895_));
  XOR2_X1   g470(.A(G301), .B(KEYINPUT88), .Z(new_n896_));
  XNOR2_X1  g471(.A(G286), .B(new_n896_), .ZN(new_n897_));
  NAND3_X1  g472(.A1(new_n894_), .A2(new_n895_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g473(.A(KEYINPUT89), .ZN(new_n899_));
  AOI21_X1  g474(.A(new_n898_), .B1(new_n899_), .B2(new_n887_), .ZN(new_n900_));
  AOI21_X1  g475(.A(new_n897_), .B1(new_n887_), .B2(KEYINPUT89), .ZN(new_n901_));
  NOR2_X1   g476(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g477(.A1(new_n893_), .A2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g478(.A(new_n875_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n904_));
  NAND3_X1  g479(.A1(new_n903_), .A2(new_n866_), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g480(.A(KEYINPUT90), .ZN(new_n906_));
  NAND2_X1  g481(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g482(.A1(new_n903_), .A2(new_n904_), .A3(KEYINPUT90), .A4(new_n866_), .ZN(new_n908_));
  NAND2_X1  g483(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  XOR2_X1   g484(.A(new_n909_), .B(KEYINPUT91), .Z(G397));
  XNOR2_X1  g485(.A(KEYINPUT92), .B(G1384), .ZN(new_n911_));
  INV_X1    g486(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g487(.A(new_n912_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n913_));
  XOR2_X1   g488(.A(KEYINPUT93), .B(G40), .Z(new_n914_));
  NAND3_X1  g489(.A1(new_n805_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  OR2_X1    g490(.A1(new_n915_), .A2(KEYINPUT94), .ZN(new_n916_));
  INV_X1    g491(.A(KEYINPUT95), .ZN(new_n917_));
  OAI211_X1 g492(.A(G40), .B(new_n912_), .C1(new_n496_), .C2(new_n499_), .ZN(new_n918_));
  OAI21_X1  g493(.A(new_n917_), .B1(new_n918_), .B2(new_n481_), .ZN(new_n919_));
  NAND2_X1  g494(.A1(new_n912_), .A2(G40), .ZN(new_n920_));
  AOI21_X1  g495(.A(new_n920_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n921_));
  AND4_X1   g496(.A1(KEYINPUT10), .A2(new_n465_), .A3(G125), .A4(G2105), .ZN(new_n922_));
  AOI21_X1  g497(.A(KEYINPUT10), .B1(new_n479_), .B2(G125), .ZN(new_n923_));
  NOR2_X1   g498(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g499(.A1(new_n921_), .A2(new_n924_), .A3(KEYINPUT95), .A4(new_n802_), .ZN(new_n925_));
  AOI22_X1  g500(.A1(new_n915_), .A2(KEYINPUT94), .B1(new_n919_), .B2(new_n925_), .ZN(new_n926_));
  AND2_X1   g501(.A1(new_n916_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g502(.A1(new_n723_), .A2(G2067), .ZN(new_n928_));
  NAND2_X1  g503(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  XOR2_X1   g504(.A(new_n929_), .B(KEYINPUT99), .Z(new_n930_));
  XNOR2_X1  g505(.A(KEYINPUT97), .B(G1996), .ZN(new_n931_));
  NOR2_X1   g506(.A1(new_n757_), .A2(new_n931_), .ZN(new_n932_));
  AND2_X1   g507(.A1(new_n927_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g508(.A(new_n931_), .ZN(new_n934_));
  NOR2_X1   g509(.A1(new_n828_), .A2(new_n934_), .ZN(new_n935_));
  OAI21_X1  g510(.A(new_n927_), .B1(new_n932_), .B2(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g511(.A(new_n936_), .B(KEYINPUT98), .ZN(new_n937_));
  INV_X1    g512(.A(new_n927_), .ZN(new_n938_));
  XNOR2_X1  g513(.A(new_n739_), .B(G1991), .ZN(new_n939_));
  NAND2_X1  g514(.A1(new_n927_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g515(.A1(G290), .A2(G1986), .ZN(new_n941_));
  NAND2_X1  g516(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  OR2_X1    g517(.A1(new_n739_), .A2(G1991), .ZN(new_n943_));
  AOI21_X1  g518(.A(new_n938_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g519(.A(new_n933_), .B1(new_n937_), .B2(new_n944_), .ZN(new_n945_));
  INV_X1    g520(.A(G2067), .ZN(new_n946_));
  NOR2_X1   g521(.A1(new_n724_), .A2(new_n946_), .ZN(new_n947_));
  OAI21_X1  g522(.A(new_n927_), .B1(new_n928_), .B2(new_n947_), .ZN(new_n948_));
  INV_X1    g523(.A(KEYINPUT96), .ZN(new_n949_));
  XNOR2_X1  g524(.A(new_n948_), .B(new_n949_), .ZN(new_n950_));
  INV_X1    g525(.A(new_n950_), .ZN(new_n951_));
  OAI21_X1  g526(.A(new_n930_), .B1(new_n945_), .B2(new_n951_), .ZN(new_n952_));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n953_));
  XNOR2_X1  g528(.A(new_n952_), .B(new_n953_), .ZN(new_n954_));
  AND2_X1   g529(.A1(G290), .A2(G1986), .ZN(new_n955_));
  OAI211_X1 g530(.A(new_n916_), .B(new_n926_), .C1(new_n941_), .C2(new_n955_), .ZN(new_n956_));
  OAI21_X1  g531(.A(new_n940_), .B1(new_n956_), .B2(KEYINPUT123), .ZN(new_n957_));
  AOI21_X1  g532(.A(new_n957_), .B1(KEYINPUT123), .B2(new_n956_), .ZN(new_n958_));
  NAND3_X1  g533(.A1(new_n958_), .A2(new_n950_), .A3(new_n937_), .ZN(new_n959_));
  XNOR2_X1  g534(.A(new_n959_), .B(KEYINPUT124), .ZN(new_n960_));
  NAND2_X1  g535(.A1(new_n925_), .A2(new_n919_), .ZN(new_n961_));
  INV_X1    g536(.A(G1981), .ZN(new_n962_));
  NAND4_X1  g537(.A1(new_n961_), .A2(G8), .A3(new_n962_), .A4(G305), .ZN(new_n963_));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n964_));
  NAND2_X1  g539(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  INV_X1    g540(.A(G8), .ZN(new_n966_));
  AOI21_X1  g541(.A(new_n966_), .B1(new_n925_), .B2(new_n919_), .ZN(new_n967_));
  NAND4_X1  g542(.A1(new_n967_), .A2(KEYINPUT101), .A3(new_n962_), .A4(G305), .ZN(new_n968_));
  NAND2_X1  g543(.A1(new_n961_), .A2(G8), .ZN(new_n969_));
  NOR2_X1   g544(.A1(G305), .A2(new_n962_), .ZN(new_n970_));
  NOR2_X1   g545(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  NAND3_X1  g546(.A1(new_n965_), .A2(new_n968_), .A3(new_n971_), .ZN(new_n972_));
  XNOR2_X1  g547(.A(KEYINPUT106), .B(G1976), .ZN(new_n973_));
  NOR2_X1   g548(.A1(new_n969_), .A2(new_n973_), .ZN(new_n974_));
  NAND2_X1  g549(.A1(new_n961_), .A2(G288), .ZN(new_n975_));
  NAND2_X1  g550(.A1(new_n975_), .A2(KEYINPUT121), .ZN(new_n976_));
  OR2_X1    g551(.A1(new_n975_), .A2(KEYINPUT121), .ZN(new_n977_));
  NAND4_X1  g552(.A1(new_n972_), .A2(new_n974_), .A3(new_n976_), .A4(new_n977_), .ZN(new_n978_));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n979_));
  INV_X1    g554(.A(G1956), .ZN(new_n980_));
  OAI211_X1 g555(.A(KEYINPUT102), .B(new_n912_), .C1(new_n496_), .C2(new_n499_), .ZN(new_n981_));
  NAND4_X1  g556(.A1(new_n981_), .A2(G40), .A3(new_n924_), .A4(new_n802_), .ZN(new_n982_));
  AOI21_X1  g557(.A(KEYINPUT102), .B1(new_n832_), .B2(new_n912_), .ZN(new_n983_));
  OAI21_X1  g558(.A(new_n980_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n984_));
  INV_X1    g559(.A(new_n913_), .ZN(new_n985_));
  NAND4_X1  g560(.A1(new_n800_), .A2(new_n804_), .A3(new_n985_), .A4(new_n914_), .ZN(new_n986_));
  OAI21_X1  g561(.A(new_n984_), .B1(G2072), .B2(new_n986_), .ZN(new_n987_));
  XNOR2_X1  g562(.A(new_n987_), .B(new_n549_), .ZN(new_n988_));
  INV_X1    g563(.A(G1348), .ZN(new_n989_));
  OAI21_X1  g564(.A(new_n989_), .B1(new_n982_), .B2(new_n983_), .ZN(new_n990_));
  OAI21_X1  g565(.A(new_n990_), .B1(G2067), .B2(new_n986_), .ZN(new_n991_));
  AND3_X1   g566(.A1(new_n991_), .A2(KEYINPUT114), .A3(new_n581_), .ZN(new_n992_));
  AOI21_X1  g567(.A(KEYINPUT114), .B1(new_n991_), .B2(new_n581_), .ZN(new_n993_));
  NOR2_X1   g568(.A1(new_n992_), .A2(new_n993_), .ZN(new_n994_));
  AND4_X1   g569(.A1(new_n800_), .A2(new_n804_), .A3(new_n985_), .A4(new_n914_), .ZN(new_n995_));
  NAND2_X1  g570(.A1(new_n995_), .A2(new_n934_), .ZN(new_n996_));
  XOR2_X1   g571(.A(KEYINPUT117), .B(G1341), .Z(new_n997_));
  NAND2_X1  g572(.A1(new_n961_), .A2(new_n997_), .ZN(new_n998_));
  AOI21_X1  g573(.A(new_n594_), .B1(new_n996_), .B2(new_n998_), .ZN(new_n999_));
  NAND2_X1  g574(.A1(new_n991_), .A2(new_n583_), .ZN(new_n1000_));
  OAI211_X1 g575(.A(new_n582_), .B(new_n990_), .C1(G2067), .C2(new_n986_), .ZN(new_n1001_));
  NAND3_X1  g576(.A1(new_n999_), .A2(new_n1000_), .A3(new_n1001_), .ZN(new_n1002_));
  AOI21_X1  g577(.A(new_n988_), .B1(new_n994_), .B2(new_n1002_), .ZN(new_n1003_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004_));
  NAND2_X1  g579(.A1(new_n987_), .A2(new_n1004_), .ZN(new_n1005_));
  OAI211_X1 g580(.A(new_n984_), .B(KEYINPUT115), .C1(G2072), .C2(new_n986_), .ZN(new_n1006_));
  AND4_X1   g581(.A1(KEYINPUT116), .A2(new_n1005_), .A3(new_n549_), .A4(new_n1006_), .ZN(new_n1007_));
  AOI21_X1  g582(.A(G299), .B1(new_n987_), .B2(new_n1004_), .ZN(new_n1008_));
  AOI21_X1  g583(.A(KEYINPUT116), .B1(new_n1008_), .B2(new_n1006_), .ZN(new_n1009_));
  NOR2_X1   g584(.A1(new_n1007_), .A2(new_n1009_), .ZN(new_n1010_));
  OAI21_X1  g585(.A(new_n979_), .B1(new_n1003_), .B2(new_n1010_), .ZN(new_n1011_));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n1012_));
  NOR2_X1   g587(.A1(new_n982_), .A2(new_n983_), .ZN(new_n1013_));
  NAND3_X1  g588(.A1(new_n1013_), .A2(KEYINPUT103), .A3(new_n808_), .ZN(new_n1014_));
  INV_X1    g589(.A(KEYINPUT103), .ZN(new_n1015_));
  INV_X1    g590(.A(KEYINPUT102), .ZN(new_n1016_));
  NAND2_X1  g591(.A1(new_n913_), .A2(new_n1016_), .ZN(new_n1017_));
  NAND4_X1  g592(.A1(new_n1017_), .A2(G160), .A3(G40), .A4(new_n981_), .ZN(new_n1018_));
  OAI21_X1  g593(.A(new_n1015_), .B1(new_n1018_), .B2(G2084), .ZN(new_n1019_));
  INV_X1    g594(.A(G1966), .ZN(new_n1020_));
  NAND2_X1  g595(.A1(new_n986_), .A2(new_n1020_), .ZN(new_n1021_));
  NAND3_X1  g596(.A1(new_n1014_), .A2(new_n1019_), .A3(new_n1021_), .ZN(new_n1022_));
  NAND2_X1  g597(.A1(G286), .A2(G8), .ZN(new_n1023_));
  XNOR2_X1  g598(.A(new_n1023_), .B(KEYINPUT104), .ZN(new_n1024_));
  NAND3_X1  g599(.A1(new_n1022_), .A2(new_n1024_), .A3(G8), .ZN(new_n1025_));
  NAND2_X1  g600(.A1(new_n1025_), .A2(new_n972_), .ZN(new_n1026_));
  AOI21_X1  g601(.A(new_n1024_), .B1(new_n1022_), .B2(G8), .ZN(new_n1027_));
  OAI21_X1  g602(.A(new_n1012_), .B1(new_n1026_), .B2(new_n1027_), .ZN(new_n1028_));
  INV_X1    g603(.A(new_n1027_), .ZN(new_n1029_));
  NAND4_X1  g604(.A1(new_n1029_), .A2(KEYINPUT105), .A3(new_n1025_), .A4(new_n972_), .ZN(new_n1030_));
  NAND2_X1  g605(.A1(new_n1028_), .A2(new_n1030_), .ZN(new_n1031_));
  INV_X1    g606(.A(new_n988_), .ZN(new_n1032_));
  AND3_X1   g607(.A1(new_n999_), .A2(new_n1001_), .A3(new_n1000_), .ZN(new_n1033_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n1034_));
  AOI22_X1  g609(.A1(new_n995_), .A2(new_n946_), .B1(new_n989_), .B2(new_n1018_), .ZN(new_n1035_));
  OAI21_X1  g610(.A(new_n1034_), .B1(new_n1035_), .B2(new_n596_), .ZN(new_n1036_));
  NAND3_X1  g611(.A1(new_n991_), .A2(KEYINPUT114), .A3(new_n581_), .ZN(new_n1037_));
  NAND2_X1  g612(.A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1038_));
  OAI21_X1  g613(.A(new_n1032_), .B1(new_n1033_), .B2(new_n1038_), .ZN(new_n1039_));
  NAND2_X1  g614(.A1(new_n1008_), .A2(new_n1006_), .ZN(new_n1040_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041_));
  NAND2_X1  g616(.A1(new_n1040_), .A2(new_n1041_), .ZN(new_n1042_));
  NAND3_X1  g617(.A1(new_n1008_), .A2(KEYINPUT116), .A3(new_n1006_), .ZN(new_n1043_));
  NAND2_X1  g618(.A1(new_n1042_), .A2(new_n1043_), .ZN(new_n1044_));
  NAND3_X1  g619(.A1(new_n1039_), .A2(new_n1044_), .A3(KEYINPUT118), .ZN(new_n1045_));
  NAND3_X1  g620(.A1(new_n1011_), .A2(new_n1031_), .A3(new_n1045_), .ZN(new_n1046_));
  OAI22_X1  g621(.A1(new_n995_), .A2(G1971), .B1(G2090), .B2(new_n1018_), .ZN(new_n1047_));
  NAND4_X1  g622(.A1(new_n1047_), .A2(KEYINPUT112), .A3(G8), .A4(G303), .ZN(new_n1048_));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049_));
  INV_X1    g624(.A(G2090), .ZN(new_n1050_));
  AOI22_X1  g625(.A1(new_n1050_), .A2(new_n1013_), .B1(new_n986_), .B2(new_n733_), .ZN(new_n1051_));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052_));
  OAI21_X1  g627(.A(new_n1049_), .B1(new_n1051_), .B2(new_n1052_), .ZN(new_n1053_));
  AOI21_X1  g628(.A(new_n966_), .B1(new_n1051_), .B2(G166), .ZN(new_n1054_));
  NAND3_X1  g629(.A1(new_n1048_), .A2(new_n1053_), .A3(new_n1054_), .ZN(new_n1055_));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n1056_));
  NAND2_X1  g631(.A1(new_n1055_), .A2(new_n1056_), .ZN(new_n1057_));
  NAND4_X1  g632(.A1(new_n1048_), .A2(new_n1053_), .A3(new_n1054_), .A4(KEYINPUT113), .ZN(new_n1058_));
  NAND2_X1  g633(.A1(new_n1057_), .A2(new_n1058_), .ZN(new_n1059_));
  AOI21_X1  g634(.A(new_n969_), .B1(new_n692_), .B2(new_n973_), .ZN(new_n1060_));
  INV_X1    g635(.A(new_n973_), .ZN(new_n1061_));
  NAND4_X1  g636(.A1(new_n967_), .A2(KEYINPUT107), .A3(G288), .A4(new_n1061_), .ZN(new_n1062_));
  NAND4_X1  g637(.A1(new_n961_), .A2(G8), .A3(G288), .A4(new_n1061_), .ZN(new_n1063_));
  INV_X1    g638(.A(KEYINPUT107), .ZN(new_n1064_));
  NAND2_X1  g639(.A1(new_n1063_), .A2(new_n1064_), .ZN(new_n1065_));
  NAND3_X1  g640(.A1(new_n1060_), .A2(new_n1062_), .A3(new_n1065_), .ZN(new_n1066_));
  XNOR2_X1  g641(.A(new_n1066_), .B(KEYINPUT108), .ZN(new_n1067_));
  XNOR2_X1  g642(.A(KEYINPUT110), .B(G1961), .ZN(new_n1068_));
  NAND2_X1  g643(.A1(new_n1018_), .A2(new_n1068_), .ZN(new_n1069_));
  INV_X1    g644(.A(new_n1069_), .ZN(new_n1070_));
  OR3_X1    g645(.A1(new_n986_), .A2(KEYINPUT109), .A3(G2078), .ZN(new_n1071_));
  OAI21_X1  g646(.A(KEYINPUT109), .B1(new_n986_), .B2(G2078), .ZN(new_n1072_));
  AOI21_X1  g647(.A(new_n1070_), .B1(new_n1071_), .B2(new_n1072_), .ZN(new_n1073_));
  NOR2_X1   g648(.A1(new_n1073_), .A2(G301), .ZN(new_n1074_));
  INV_X1    g649(.A(new_n1074_), .ZN(new_n1075_));
  AOI211_X1 g650(.A(G171), .B(new_n1070_), .C1(new_n1071_), .C2(new_n1072_), .ZN(new_n1076_));
  INV_X1    g651(.A(new_n1076_), .ZN(new_n1077_));
  AOI21_X1  g652(.A(KEYINPUT111), .B1(new_n1075_), .B2(new_n1077_), .ZN(new_n1078_));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n1079_));
  NOR3_X1   g654(.A1(new_n1074_), .A2(new_n1076_), .A3(new_n1079_), .ZN(new_n1080_));
  OAI211_X1 g655(.A(new_n1059_), .B(new_n1067_), .C1(new_n1078_), .C2(new_n1080_), .ZN(new_n1081_));
  OAI21_X1  g656(.A(new_n978_), .B1(new_n1046_), .B2(new_n1081_), .ZN(new_n1082_));
  NOR3_X1   g657(.A1(new_n969_), .A2(G1981), .A3(G305), .ZN(new_n1083_));
  INV_X1    g658(.A(new_n972_), .ZN(new_n1084_));
  NOR4_X1   g659(.A1(new_n1084_), .A2(new_n966_), .A3(G303), .A4(new_n1051_), .ZN(new_n1085_));
  AOI21_X1  g660(.A(new_n1083_), .B1(new_n1085_), .B2(new_n1067_), .ZN(new_n1086_));
  OAI21_X1  g661(.A(KEYINPUT119), .B1(new_n1073_), .B2(G301), .ZN(new_n1087_));
  AND2_X1   g662(.A1(new_n1087_), .A2(new_n1066_), .ZN(new_n1088_));
  NOR2_X1   g663(.A1(new_n1026_), .A2(new_n1027_), .ZN(new_n1089_));
  OR3_X1    g664(.A1(new_n1073_), .A2(KEYINPUT119), .A3(G301), .ZN(new_n1090_));
  NAND4_X1  g665(.A1(new_n1059_), .A2(new_n1088_), .A3(new_n1089_), .A4(new_n1090_), .ZN(new_n1091_));
  NOR2_X1   g666(.A1(new_n1084_), .A2(new_n1025_), .ZN(new_n1092_));
  NAND3_X1  g667(.A1(new_n1059_), .A2(new_n1067_), .A3(new_n1092_), .ZN(new_n1093_));
  NAND3_X1  g668(.A1(new_n1086_), .A2(new_n1091_), .A3(new_n1093_), .ZN(new_n1094_));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095_));
  NAND2_X1  g670(.A1(new_n1094_), .A2(new_n1095_), .ZN(new_n1096_));
  NAND4_X1  g671(.A1(new_n1086_), .A2(new_n1091_), .A3(new_n1093_), .A4(KEYINPUT120), .ZN(new_n1097_));
  AOI21_X1  g672(.A(new_n1082_), .B1(new_n1096_), .B2(new_n1097_), .ZN(new_n1098_));
  OAI21_X1  g673(.A(new_n960_), .B1(new_n1098_), .B2(KEYINPUT122), .ZN(new_n1099_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100_));
  AOI211_X1 g675(.A(new_n1100_), .B(new_n1082_), .C1(new_n1096_), .C2(new_n1097_), .ZN(new_n1101_));
  OAI21_X1  g676(.A(new_n954_), .B1(new_n1099_), .B2(new_n1101_), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g677(.A1(new_n669_), .A2(new_n632_), .A3(new_n670_), .ZN(new_n1104_));
  AOI21_X1  g678(.A(new_n459_), .B1(new_n1104_), .B2(KEYINPUT126), .ZN(new_n1105_));
  OAI21_X1  g679(.A(new_n1105_), .B1(KEYINPUT126), .B2(new_n1104_), .ZN(new_n1106_));
  AOI21_X1  g680(.A(new_n1106_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n1107_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n1108_));
  INV_X1    g682(.A(G227), .ZN(new_n1109_));
  AND3_X1   g683(.A1(new_n869_), .A2(new_n1108_), .A3(new_n1109_), .ZN(new_n1110_));
  AOI21_X1  g684(.A(new_n1108_), .B1(new_n869_), .B2(new_n1109_), .ZN(new_n1111_));
  OAI21_X1  g685(.A(new_n1107_), .B1(new_n1110_), .B2(new_n1111_), .ZN(G225));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n1113_));
  NAND2_X1  g687(.A1(G225), .A2(new_n1113_), .ZN(new_n1114_));
  OAI211_X1 g688(.A(new_n1107_), .B(KEYINPUT127), .C1(new_n1110_), .C2(new_n1111_), .ZN(new_n1115_));
  NAND2_X1  g689(.A1(new_n1114_), .A2(new_n1115_), .ZN(G308));
endmodule


