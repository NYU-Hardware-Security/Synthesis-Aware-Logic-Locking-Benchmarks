//Secret key is'0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_c5315" written by ABC on Mon Oct 31 10:37:46 2022

module locked_c5315 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G4, G11, G14, G17,
    G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52,
    G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86,
    G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149,
    G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185,
    G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225,
    G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265,
    G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308,
    G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358,
    G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435,
    G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552,
    G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358,
    G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088,
    G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G4,
    G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43,
    G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81,
    G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145,
    G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179,
    G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217,
    G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257,
    G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302,
    G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348,
    G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411,
    G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545,
    G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174,
    G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087,
    G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_n384_, new_n386_, new_n396_, new_n404_, new_n406_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n415_, new_n416_, new_n418_,
    new_n419_, new_n421_, new_n422_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1107_, new_n1108_, new_n1110_, new_n1111_, new_n1112_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1122_, new_n1123_, new_n1124_, new_n1126_, new_n1127_,
    new_n1129_, new_n1130_, new_n1131_, new_n1133_, new_n1134_, new_n1135_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_;
  BUF_X1    g0000(.A(G141), .Z(G144));
  BUF_X1    g0001(.A(G293), .Z(G298));
  BUF_X1    g0002(.A(G3173), .Z(G973));
  INV_X1    g0003(.A(G545), .ZN(G594));
  INV_X1    g0004(.A(G348), .ZN(G599));
  INV_X1    g0005(.A(G366), .ZN(G600));
  INV_X1    g0006(.A(G552), .ZN(G849));
  INV_X1    g0007(.A(G562), .ZN(G850));
  NOR2_X1   g0008(.A1(G849), .A2(G850), .ZN(G601));
  INV_X1    g0009(.A(G549), .ZN(G602));
  INV_X1    g0010(.A(G545), .ZN(G603));
  INV_X1    g0011(.A(G545), .ZN(G604));
  XNOR2_X1  g0012(.A(KEYINPUT0), .B(G338), .ZN(G611));
  INV_X1    g0013(.A(G358), .ZN(G612));
  AND2_X1   g0014(.A1(G141), .A2(G145), .ZN(G810));
  INV_X1    g0015(.A(G245), .ZN(G848));
  INV_X1    g0016(.A(G559), .ZN(G851));
  AND2_X1   g0017(.A1(G1), .A2(G373), .ZN(G634));
  INV_X1    g0018(.A(G136), .ZN(new_n384_));
  NOR2_X1   g0019(.A1(new_n384_), .A2(G3173), .ZN(G815));
  INV_X1    g0020(.A(G2824), .ZN(new_n386_));
  NAND2_X1  g0021(.A1(new_n386_), .A2(G27), .ZN(G845));
  NAND2_X1  g0022(.A1(G386), .A2(G556), .ZN(G847));
  BUF_X1    g0023(.A(G137), .Z(G926));
  BUF_X1    g0024(.A(G141), .Z(G923));
  BUF_X1    g0025(.A(G1), .Z(G921));
  XNOR2_X1  g0026(.A(KEYINPUT1), .B(G549), .ZN(G892));
  BUF_X1    g0027(.A(G299), .Z(G887));
  INV_X1    g0028(.A(G549), .ZN(G606));
  NAND2_X1  g0029(.A1(G27), .A2(G31), .ZN(G809));
  INV_X1    g0030(.A(G809), .ZN(new_n396_));
  NAND2_X1  g0031(.A1(new_n396_), .A2(G140), .ZN(G656));
  BUF_X1    g0032(.A(G1), .Z(G993));
  BUF_X1    g0033(.A(G1), .Z(G978));
  BUF_X1    g0034(.A(G1), .Z(G949));
  BUF_X1    g0035(.A(G1), .Z(G939));
  BUF_X1    g0036(.A(G299), .Z(G889));
  INV_X1    g0037(.A(G299), .ZN(G593));
  MUX2_X1   g0038(.A(G86), .B(G87), .S(G2358), .Z(new_n404_));
  NAND2_X1  g0039(.A1(new_n404_), .A2(new_n396_), .ZN(G636));
  MUX2_X1   g0040(.A(G88), .B(G34), .S(G2358), .Z(new_n406_));
  NAND2_X1  g0041(.A1(new_n406_), .A2(new_n396_), .ZN(G704));
  NAND2_X1  g0042(.A1(new_n406_), .A2(new_n396_), .ZN(G717));
  NAND2_X1  g0043(.A1(new_n396_), .A2(G83), .ZN(G820));
  INV_X1    g0044(.A(G141), .ZN(new_n410_));
  XOR2_X1   g0045(.A(KEYINPUT2), .B(G2358), .Z(new_n411_));
  NAND2_X1  g0046(.A1(new_n411_), .A2(G24), .ZN(new_n412_));
  AOI21_X1  g0047(.A(G809), .B1(G25), .B2(G2358), .ZN(new_n413_));
  AOI21_X1  g0048(.A(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(G639));
  NAND2_X1  g0049(.A1(new_n411_), .A2(G26), .ZN(new_n415_));
  AOI21_X1  g0050(.A(G809), .B1(G81), .B2(G2358), .ZN(new_n416_));
  AOI21_X1  g0051(.A(new_n410_), .B1(new_n415_), .B2(new_n416_), .ZN(G673));
  NAND2_X1  g0052(.A1(new_n411_), .A2(G79), .ZN(new_n418_));
  AOI21_X1  g0053(.A(G809), .B1(G23), .B2(G2358), .ZN(new_n419_));
  AOI21_X1  g0054(.A(new_n410_), .B1(new_n418_), .B2(new_n419_), .ZN(G707));
  NAND2_X1  g0055(.A1(new_n411_), .A2(G82), .ZN(new_n421_));
  AOI21_X1  g0056(.A(G809), .B1(G80), .B2(G2358), .ZN(new_n422_));
  AOI21_X1  g0057(.A(new_n410_), .B1(new_n421_), .B2(new_n422_), .ZN(G715));
  INV_X1    g0058(.A(G479), .ZN(new_n424_));
  INV_X1    g0059(.A(G308), .ZN(new_n425_));
  NOR2_X1   g0060(.A1(new_n425_), .A2(G242), .ZN(new_n426_));
  NOR2_X1   g0061(.A1(G254), .A2(G308), .ZN(new_n427_));
  OAI21_X1  g0062(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g0063(.A(G251), .ZN(new_n429_));
  INV_X1    g0064(.A(G248), .ZN(new_n430_));
  MUX2_X1   g0065(.A(new_n429_), .B(new_n430_), .S(G308), .Z(new_n431_));
  OAI21_X1  g0066(.A(new_n428_), .B1(new_n431_), .B2(new_n424_), .ZN(new_n432_));
  INV_X1    g0067(.A(G490), .ZN(new_n433_));
  INV_X1    g0068(.A(G316), .ZN(new_n434_));
  NOR2_X1   g0069(.A1(new_n434_), .A2(G242), .ZN(new_n435_));
  NOR2_X1   g0070(.A1(G254), .A2(G316), .ZN(new_n436_));
  OAI21_X1  g0071(.A(new_n433_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  MUX2_X1   g0072(.A(new_n429_), .B(new_n430_), .S(G316), .Z(new_n438_));
  OAI21_X1  g0073(.A(new_n437_), .B1(new_n438_), .B2(new_n433_), .ZN(new_n439_));
  NAND2_X1  g0074(.A1(G242), .A2(G293), .ZN(new_n440_));
  INV_X1    g0075(.A(G254), .ZN(new_n441_));
  OAI21_X1  g0076(.A(new_n440_), .B1(new_n441_), .B2(G293), .ZN(new_n442_));
  INV_X1    g0077(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g0078(.A1(G248), .A2(G302), .ZN(new_n444_));
  OAI21_X1  g0079(.A(new_n444_), .B1(new_n429_), .B2(G302), .ZN(new_n445_));
  AND2_X1   g0080(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g0081(.A1(G248), .A2(G361), .ZN(new_n447_));
  OAI21_X1  g0082(.A(new_n447_), .B1(new_n429_), .B2(G361), .ZN(new_n448_));
  AND4_X1   g0083(.A1(new_n432_), .A2(new_n439_), .A3(new_n446_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g0084(.A(G523), .ZN(new_n450_));
  XOR2_X1   g0085(.A(KEYINPUT3), .B(G341), .Z(new_n451_));
  INV_X1    g0086(.A(new_n451_), .ZN(new_n452_));
  OAI221_X1 g0087(.A(new_n450_), .B1(G341), .B2(G3548), .C1(new_n452_), .C2(G3546), .ZN(new_n453_));
  INV_X1    g0088(.A(G3550), .ZN(new_n454_));
  INV_X1    g0089(.A(G3552), .ZN(new_n455_));
  AOI22_X1  g0090(.A1(new_n452_), .A2(new_n454_), .B1(G341), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g0091(.A(new_n453_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g0092(.A(G324), .ZN(new_n458_));
  NOR2_X1   g0093(.A1(new_n458_), .A2(G3552), .ZN(new_n459_));
  NOR2_X1   g0094(.A1(G324), .A2(G3550), .ZN(new_n460_));
  OAI21_X1  g0095(.A(G503), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g0096(.A(G3548), .ZN(new_n462_));
  INV_X1    g0097(.A(G3546), .ZN(new_n463_));
  MUX2_X1   g0098(.A(new_n462_), .B(new_n463_), .S(G324), .Z(new_n464_));
  OAI21_X1  g0099(.A(new_n461_), .B1(new_n464_), .B2(G503), .ZN(new_n465_));
  NAND2_X1  g0100(.A1(new_n455_), .A2(G514), .ZN(new_n466_));
  OAI21_X1  g0101(.A(new_n466_), .B1(G514), .B2(new_n463_), .ZN(new_n467_));
  INV_X1    g0102(.A(G351), .ZN(new_n468_));
  NOR2_X1   g0103(.A1(new_n468_), .A2(G3552), .ZN(new_n469_));
  NOR2_X1   g0104(.A1(G351), .A2(G3550), .ZN(new_n470_));
  OAI21_X1  g0105(.A(G534), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  MUX2_X1   g0106(.A(new_n462_), .B(new_n463_), .S(G351), .Z(new_n472_));
  OAI21_X1  g0107(.A(new_n471_), .B1(new_n472_), .B2(G534), .ZN(new_n473_));
  NAND4_X1  g0108(.A1(new_n457_), .A2(new_n465_), .A3(new_n467_), .A4(new_n473_), .ZN(new_n474_));
  OAI21_X1  g0109(.A(new_n449_), .B1(new_n474_), .B2(KEYINPUT4), .ZN(new_n475_));
  AOI21_X1  g0110(.A(new_n475_), .B1(KEYINPUT4), .B2(new_n474_), .ZN(G598));
  NAND3_X1  g0111(.A1(new_n455_), .A2(G218), .A3(G468), .ZN(new_n477_));
  XOR2_X1   g0112(.A(new_n477_), .B(KEYINPUT5), .Z(new_n478_));
  INV_X1    g0113(.A(G218), .ZN(new_n479_));
  NAND3_X1  g0114(.A1(new_n479_), .A2(new_n454_), .A3(G468), .ZN(new_n480_));
  MUX2_X1   g0115(.A(new_n462_), .B(new_n463_), .S(G218), .Z(new_n481_));
  OAI211_X1 g0116(.A(new_n478_), .B(new_n480_), .C1(G468), .C2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g0117(.A(new_n482_), .B(KEYINPUT6), .Z(new_n483_));
  INV_X1    g0118(.A(G265), .ZN(new_n484_));
  NOR2_X1   g0119(.A1(new_n484_), .A2(G3552), .ZN(new_n485_));
  NOR2_X1   g0120(.A1(G265), .A2(G3550), .ZN(new_n486_));
  OAI21_X1  g0121(.A(G400), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  MUX2_X1   g0122(.A(new_n462_), .B(new_n463_), .S(G265), .Z(new_n488_));
  OAI21_X1  g0123(.A(new_n487_), .B1(new_n488_), .B2(G400), .ZN(new_n489_));
  INV_X1    g0124(.A(G257), .ZN(new_n490_));
  NOR2_X1   g0125(.A1(new_n490_), .A2(G3552), .ZN(new_n491_));
  NOR2_X1   g0126(.A1(G257), .A2(G3550), .ZN(new_n492_));
  OAI21_X1  g0127(.A(G389), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  MUX2_X1   g0128(.A(new_n462_), .B(new_n463_), .S(G257), .Z(new_n494_));
  OAI21_X1  g0129(.A(new_n493_), .B1(new_n494_), .B2(G389), .ZN(new_n495_));
  INV_X1    g0130(.A(G210), .ZN(new_n496_));
  NOR2_X1   g0131(.A1(new_n496_), .A2(G3552), .ZN(new_n497_));
  NOR2_X1   g0132(.A1(G210), .A2(G3550), .ZN(new_n498_));
  OAI21_X1  g0133(.A(G457), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  MUX2_X1   g0134(.A(new_n462_), .B(new_n463_), .S(G210), .Z(new_n500_));
  OAI21_X1  g0135(.A(new_n499_), .B1(new_n500_), .B2(G457), .ZN(new_n501_));
  AND3_X1   g0136(.A1(new_n489_), .A2(new_n495_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g0137(.A1(new_n455_), .A2(G234), .A3(G435), .ZN(new_n503_));
  XNOR2_X1  g0138(.A(new_n503_), .B(KEYINPUT7), .ZN(new_n504_));
  INV_X1    g0139(.A(G234), .ZN(new_n505_));
  NAND3_X1  g0140(.A1(new_n505_), .A2(new_n454_), .A3(G435), .ZN(new_n506_));
  MUX2_X1   g0141(.A(new_n462_), .B(new_n463_), .S(G234), .Z(new_n507_));
  OAI211_X1 g0142(.A(new_n504_), .B(new_n506_), .C1(G435), .C2(new_n507_), .ZN(new_n508_));
  INV_X1    g0143(.A(G422), .ZN(new_n509_));
  INV_X1    g0144(.A(G226), .ZN(new_n510_));
  NAND2_X1  g0145(.A1(new_n510_), .A2(new_n454_), .ZN(new_n511_));
  NAND2_X1  g0146(.A1(new_n455_), .A2(G226), .ZN(new_n512_));
  AOI21_X1  g0147(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g0148(.A1(new_n510_), .A2(G3548), .ZN(new_n514_));
  NAND2_X1  g0149(.A1(G226), .A2(G3546), .ZN(new_n515_));
  AOI21_X1  g0150(.A(G422), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g0151(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g0152(.A(G411), .ZN(new_n518_));
  INV_X1    g0153(.A(G273), .ZN(new_n519_));
  NAND2_X1  g0154(.A1(new_n519_), .A2(new_n454_), .ZN(new_n520_));
  NAND2_X1  g0155(.A1(new_n455_), .A2(G273), .ZN(new_n521_));
  AOI21_X1  g0156(.A(new_n518_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g0157(.A1(new_n519_), .A2(G3548), .ZN(new_n523_));
  NAND2_X1  g0158(.A1(G273), .A2(G3546), .ZN(new_n524_));
  AOI21_X1  g0159(.A(G411), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g0160(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g0161(.A(G206), .ZN(new_n527_));
  NAND2_X1  g0162(.A1(new_n527_), .A2(new_n441_), .ZN(new_n528_));
  INV_X1    g0163(.A(G242), .ZN(new_n529_));
  NAND2_X1  g0164(.A1(new_n529_), .A2(G206), .ZN(new_n530_));
  AOI21_X1  g0165(.A(G446), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g0166(.A(G446), .ZN(new_n532_));
  NAND2_X1  g0167(.A1(new_n527_), .A2(G251), .ZN(new_n533_));
  NAND2_X1  g0168(.A1(G206), .A2(G248), .ZN(new_n534_));
  AOI21_X1  g0169(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g0170(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g0171(.A(G374), .ZN(new_n537_));
  INV_X1    g0172(.A(G281), .ZN(new_n538_));
  NAND2_X1  g0173(.A1(new_n538_), .A2(new_n454_), .ZN(new_n539_));
  NAND2_X1  g0174(.A1(new_n455_), .A2(G281), .ZN(new_n540_));
  AOI21_X1  g0175(.A(new_n537_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g0176(.A1(new_n538_), .A2(G3548), .ZN(new_n542_));
  NAND2_X1  g0177(.A1(G281), .A2(G3546), .ZN(new_n543_));
  AOI21_X1  g0178(.A(G374), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g0179(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NOR4_X1   g0180(.A1(new_n517_), .A2(new_n526_), .A3(new_n536_), .A4(new_n545_), .ZN(new_n546_));
  AND4_X1   g0181(.A1(new_n483_), .A2(new_n502_), .A3(new_n508_), .A4(new_n546_), .ZN(G610));
  INV_X1    g0182(.A(G335), .ZN(new_n548_));
  NAND2_X1  g0183(.A1(new_n548_), .A2(G265), .ZN(new_n549_));
  NAND2_X1  g0184(.A1(G272), .A2(G335), .ZN(new_n550_));
  AND2_X1   g0185(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g0186(.A(G400), .ZN(new_n552_));
  NAND2_X1  g0187(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g0188(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g0189(.A1(new_n551_), .A2(new_n552_), .ZN(new_n555_));
  NOR2_X1   g0190(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g0191(.A1(new_n548_), .A2(G257), .ZN(new_n557_));
  NAND2_X1  g0192(.A1(G264), .A2(G335), .ZN(new_n558_));
  NAND2_X1  g0193(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g0194(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g0195(.A(G389), .ZN(new_n561_));
  NAND2_X1  g0196(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g0197(.A1(new_n559_), .A2(G389), .ZN(new_n563_));
  NAND2_X1  g0198(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g0199(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g0200(.A1(new_n556_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g0201(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g0202(.A1(new_n505_), .A2(G335), .ZN(new_n568_));
  AOI21_X1  g0203(.A(new_n568_), .B1(G241), .B2(G335), .ZN(new_n569_));
  INV_X1    g0204(.A(G435), .ZN(new_n570_));
  NOR2_X1   g0205(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g0206(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g0207(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  NAND2_X1  g0208(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g0209(.A(new_n574_), .ZN(new_n575_));
  AND2_X1   g0210(.A1(G288), .A2(G335), .ZN(new_n576_));
  AOI21_X1  g0211(.A(new_n576_), .B1(G281), .B2(new_n548_), .ZN(new_n577_));
  NOR2_X1   g0212(.A1(new_n577_), .A2(new_n537_), .ZN(new_n578_));
  INV_X1    g0213(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g0214(.A1(new_n548_), .A2(G273), .ZN(new_n580_));
  NAND2_X1  g0215(.A1(G280), .A2(G335), .ZN(new_n581_));
  AND2_X1   g0216(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g0217(.A1(new_n582_), .A2(G411), .ZN(new_n583_));
  NAND2_X1  g0218(.A1(new_n580_), .A2(new_n581_), .ZN(new_n584_));
  NAND2_X1  g0219(.A1(new_n584_), .A2(new_n518_), .ZN(new_n585_));
  NAND2_X1  g0220(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g0221(.A1(new_n577_), .A2(new_n537_), .ZN(new_n587_));
  NAND3_X1  g0222(.A1(new_n579_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g0223(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g0224(.A1(new_n567_), .A2(new_n575_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g0225(.A1(new_n548_), .A2(G226), .ZN(new_n591_));
  NAND2_X1  g0226(.A1(G233), .A2(G335), .ZN(new_n592_));
  AND2_X1   g0227(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g0228(.A1(new_n593_), .A2(new_n509_), .ZN(new_n594_));
  INV_X1    g0229(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g0230(.A1(new_n593_), .A2(new_n509_), .ZN(new_n596_));
  NAND2_X1  g0231(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g0232(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g0233(.A1(new_n527_), .A2(G335), .ZN(new_n599_));
  AOI21_X1  g0234(.A(new_n599_), .B1(G209), .B2(G335), .ZN(new_n600_));
  NAND2_X1  g0235(.A1(new_n600_), .A2(new_n532_), .ZN(new_n601_));
  INV_X1    g0236(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g0237(.A1(new_n600_), .A2(new_n532_), .ZN(new_n603_));
  NOR2_X1   g0238(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g0239(.A1(G217), .A2(G335), .ZN(new_n605_));
  OAI21_X1  g0240(.A(new_n605_), .B1(new_n496_), .B2(G335), .ZN(new_n606_));
  OR2_X1    g0241(.A1(new_n606_), .A2(G457), .ZN(new_n607_));
  NAND2_X1  g0242(.A1(new_n606_), .A2(G457), .ZN(new_n608_));
  NAND2_X1  g0243(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g0244(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g0245(.A1(G225), .A2(G335), .ZN(new_n611_));
  OAI21_X1  g0246(.A(new_n611_), .B1(new_n479_), .B2(G335), .ZN(new_n612_));
  INV_X1    g0247(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g0248(.A(G468), .ZN(new_n614_));
  NAND2_X1  g0249(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g0250(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g0251(.A1(new_n612_), .A2(G468), .ZN(new_n617_));
  INV_X1    g0252(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g0253(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g0254(.A1(new_n598_), .A2(new_n604_), .A3(new_n610_), .A4(new_n619_), .ZN(new_n620_));
  NOR2_X1   g0255(.A1(new_n590_), .A2(new_n620_), .ZN(G588));
  INV_X1    g0256(.A(KEYINPUT10), .ZN(new_n622_));
  NAND2_X1  g0257(.A1(G332), .A2(G358), .ZN(new_n623_));
  INV_X1    g0258(.A(G534), .ZN(new_n624_));
  OAI211_X1 g0259(.A(new_n623_), .B(new_n624_), .C1(G332), .C2(new_n468_), .ZN(new_n625_));
  INV_X1    g0260(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g0261(.A(G332), .ZN(new_n627_));
  NAND2_X1  g0262(.A1(new_n627_), .A2(G351), .ZN(new_n628_));
  AOI21_X1  g0263(.A(new_n624_), .B1(new_n628_), .B2(new_n623_), .ZN(new_n629_));
  OAI21_X1  g0264(.A(new_n622_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g0265(.A(new_n623_), .B1(new_n468_), .B2(G332), .ZN(new_n631_));
  NAND2_X1  g0266(.A1(new_n631_), .A2(G534), .ZN(new_n632_));
  NAND3_X1  g0267(.A1(new_n632_), .A2(KEYINPUT10), .A3(new_n625_), .ZN(new_n633_));
  NAND2_X1  g0268(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g0269(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g0270(.A1(G332), .A2(G348), .ZN(new_n636_));
  INV_X1    g0271(.A(G341), .ZN(new_n637_));
  OAI21_X1  g0272(.A(new_n636_), .B1(new_n637_), .B2(G332), .ZN(new_n638_));
  INV_X1    g0273(.A(new_n638_), .ZN(new_n639_));
  NOR2_X1   g0274(.A1(new_n639_), .A2(new_n450_), .ZN(new_n640_));
  INV_X1    g0275(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g0276(.A1(G611), .A2(G332), .ZN(new_n642_));
  NAND3_X1  g0277(.A1(new_n642_), .A2(KEYINPUT9), .A3(G514), .ZN(new_n643_));
  NAND2_X1  g0278(.A1(new_n639_), .A2(new_n450_), .ZN(new_n644_));
  XOR2_X1   g0279(.A(KEYINPUT9), .B(G514), .Z(new_n645_));
  NAND3_X1  g0280(.A1(new_n645_), .A2(G332), .A3(G611), .ZN(new_n646_));
  NAND4_X1  g0281(.A1(new_n641_), .A2(new_n643_), .A3(new_n644_), .A4(new_n646_), .ZN(new_n647_));
  NOR2_X1   g0282(.A1(new_n635_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g0283(.A1(G331), .A2(G332), .ZN(new_n649_));
  OAI21_X1  g0284(.A(new_n649_), .B1(new_n458_), .B2(G332), .ZN(new_n650_));
  INV_X1    g0285(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g0286(.A(G503), .ZN(new_n652_));
  NAND2_X1  g0287(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g0288(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g0289(.A1(new_n651_), .A2(new_n652_), .ZN(new_n655_));
  NOR2_X1   g0290(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g0291(.A1(G332), .A2(G366), .ZN(new_n657_));
  INV_X1    g0292(.A(G361), .ZN(new_n658_));
  OAI21_X1  g0293(.A(new_n657_), .B1(new_n658_), .B2(G332), .ZN(new_n659_));
  INV_X1    g0294(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g0295(.A1(new_n648_), .A2(new_n656_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0296(.A1(new_n627_), .A2(G316), .ZN(new_n662_));
  NAND2_X1  g0297(.A1(G323), .A2(G332), .ZN(new_n663_));
  NAND2_X1  g0298(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g0299(.A1(new_n664_), .A2(G490), .ZN(new_n665_));
  NAND2_X1  g0300(.A1(G315), .A2(G332), .ZN(new_n666_));
  OAI21_X1  g0301(.A(new_n666_), .B1(new_n425_), .B2(G332), .ZN(new_n667_));
  NAND2_X1  g0302(.A1(new_n667_), .A2(G479), .ZN(new_n668_));
  NAND2_X1  g0303(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g0304(.A(new_n667_), .ZN(new_n670_));
  NAND2_X1  g0305(.A1(new_n670_), .A2(new_n424_), .ZN(new_n671_));
  AND2_X1   g0306(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g0307(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g0308(.A1(G307), .A2(G332), .ZN(new_n674_));
  INV_X1    g0309(.A(G302), .ZN(new_n675_));
  OAI21_X1  g0310(.A(new_n674_), .B1(new_n675_), .B2(G332), .ZN(new_n676_));
  INV_X1    g0311(.A(new_n676_), .ZN(new_n677_));
  INV_X1    g0312(.A(new_n664_), .ZN(new_n678_));
  NAND2_X1  g0313(.A1(new_n678_), .A2(new_n433_), .ZN(new_n679_));
  INV_X1    g0314(.A(new_n679_), .ZN(new_n680_));
  INV_X1    g0315(.A(new_n671_), .ZN(new_n681_));
  OAI21_X1  g0316(.A(new_n668_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g0317(.A1(G299), .A2(G332), .ZN(new_n683_));
  XNOR2_X1  g0318(.A(KEYINPUT8), .B(G293), .ZN(new_n684_));
  OAI21_X1  g0319(.A(new_n683_), .B1(new_n684_), .B2(G332), .ZN(new_n685_));
  INV_X1    g0320(.A(new_n685_), .ZN(new_n686_));
  NAND4_X1  g0321(.A1(new_n673_), .A2(new_n677_), .A3(new_n682_), .A4(new_n686_), .ZN(new_n687_));
  NOR2_X1   g0322(.A1(new_n661_), .A2(new_n687_), .ZN(G615));
  NAND2_X1  g0323(.A1(new_n627_), .A2(G361), .ZN(new_n689_));
  NAND3_X1  g0324(.A1(new_n689_), .A2(KEYINPUT11), .A3(new_n657_), .ZN(new_n690_));
  INV_X1    g0325(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g0326(.A(KEYINPUT11), .B1(new_n689_), .B2(new_n657_), .ZN(new_n692_));
  NOR2_X1   g0327(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g0328(.A(new_n693_), .ZN(new_n694_));
  NAND2_X1  g0329(.A1(new_n648_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g0330(.A(new_n656_), .ZN(new_n696_));
  NOR2_X1   g0331(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g0332(.A(new_n697_), .ZN(new_n698_));
  NOR2_X1   g0333(.A1(new_n698_), .A2(new_n687_), .ZN(G626));
  XOR2_X1   g0334(.A(G588), .B(KEYINPUT12), .Z(G632));
  XNOR2_X1  g0335(.A(G308), .B(G316), .ZN(new_n701_));
  XNOR2_X1  g0336(.A(new_n701_), .B(G293), .ZN(new_n702_));
  XNOR2_X1  g0337(.A(new_n702_), .B(G302), .ZN(new_n703_));
  XOR2_X1   g0338(.A(G341), .B(G351), .Z(new_n704_));
  XNOR2_X1  g0339(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g0340(.A(G361), .B(G369), .ZN(new_n706_));
  XNOR2_X1  g0341(.A(new_n706_), .B(G324), .ZN(new_n707_));
  XNOR2_X1  g0342(.A(new_n705_), .B(new_n707_), .ZN(G1002));
  XNOR2_X1  g0343(.A(G218), .B(G226), .ZN(new_n709_));
  XNOR2_X1  g0344(.A(new_n709_), .B(G206), .ZN(new_n710_));
  XNOR2_X1  g0345(.A(new_n710_), .B(new_n496_), .ZN(new_n711_));
  XOR2_X1   g0346(.A(G265), .B(G273), .Z(new_n712_));
  XNOR2_X1  g0347(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  XOR2_X1   g0348(.A(G234), .B(G257), .Z(new_n714_));
  INV_X1    g0349(.A(new_n714_), .ZN(new_n715_));
  XOR2_X1   g0350(.A(G281), .B(G289), .Z(new_n716_));
  AOI21_X1  g0351(.A(KEYINPUT13), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g0352(.A(new_n717_), .B1(new_n716_), .B2(new_n715_), .ZN(new_n718_));
  XNOR2_X1  g0353(.A(new_n713_), .B(new_n718_), .ZN(G1004));
  INV_X1    g0354(.A(new_n603_), .ZN(new_n720_));
  NAND2_X1  g0355(.A1(new_n619_), .A2(new_n594_), .ZN(new_n721_));
  XNOR2_X1  g0356(.A(new_n617_), .B(KEYINPUT14), .ZN(new_n722_));
  NAND3_X1  g0357(.A1(new_n721_), .A2(new_n610_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g0358(.A1(new_n723_), .A2(new_n607_), .ZN(new_n724_));
  INV_X1    g0359(.A(new_n556_), .ZN(new_n725_));
  NOR2_X1   g0360(.A1(new_n582_), .A2(new_n518_), .ZN(new_n726_));
  INV_X1    g0361(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g0362(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g0363(.A1(new_n586_), .A2(new_n553_), .A3(new_n578_), .ZN(new_n729_));
  INV_X1    g0364(.A(new_n555_), .ZN(new_n730_));
  NAND2_X1  g0365(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g0366(.A(new_n562_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g0367(.A1(new_n732_), .A2(new_n572_), .A3(new_n563_), .ZN(new_n733_));
  NAND2_X1  g0368(.A1(new_n733_), .A2(new_n573_), .ZN(new_n734_));
  OAI221_X1 g0369(.A(new_n720_), .B1(new_n602_), .B2(new_n724_), .C1(new_n734_), .C2(new_n620_), .ZN(G591));
  NOR2_X1   g0370(.A1(new_n685_), .A2(new_n676_), .ZN(new_n736_));
  OAI211_X1 g0371(.A(new_n641_), .B(new_n632_), .C1(new_n635_), .C2(new_n694_), .ZN(new_n737_));
  NAND2_X1  g0372(.A1(new_n643_), .A2(new_n646_), .ZN(new_n738_));
  INV_X1    g0373(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g0374(.A1(new_n737_), .A2(new_n644_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g0375(.A1(new_n642_), .A2(G514), .ZN(new_n741_));
  NAND2_X1  g0376(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g0377(.A(new_n655_), .B1(new_n742_), .B2(new_n653_), .ZN(new_n743_));
  OAI211_X1 g0378(.A(new_n736_), .B(new_n673_), .C1(new_n743_), .C2(new_n687_), .ZN(G618));
  OAI221_X1 g0379(.A(new_n720_), .B1(new_n602_), .B2(new_n724_), .C1(new_n734_), .C2(new_n620_), .ZN(G621));
  OAI211_X1 g0380(.A(new_n736_), .B(new_n673_), .C1(new_n743_), .C2(new_n687_), .ZN(G629));
  INV_X1    g0381(.A(G54), .ZN(new_n747_));
  NAND2_X1  g0382(.A1(new_n660_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g0383(.A1(new_n659_), .A2(G54), .ZN(new_n749_));
  NAND2_X1  g0384(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g0385(.A1(new_n750_), .A2(G4091), .ZN(new_n751_));
  INV_X1    g0386(.A(new_n448_), .ZN(new_n752_));
  INV_X1    g0387(.A(G4091), .ZN(new_n753_));
  NAND2_X1  g0388(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g0389(.A(G4092), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g0390(.A(G4092), .ZN(new_n756_));
  NOR2_X1   g0391(.A1(new_n756_), .A2(G4091), .ZN(new_n757_));
  AOI21_X1  g0392(.A(new_n755_), .B1(G131), .B2(new_n757_), .ZN(G822));
  NOR3_X1   g0393(.A1(new_n473_), .A2(G4091), .A3(G4092), .ZN(new_n759_));
  AND2_X1   g0394(.A1(new_n634_), .A2(new_n748_), .ZN(new_n760_));
  NOR2_X1   g0395(.A1(new_n634_), .A2(new_n748_), .ZN(new_n761_));
  NOR2_X1   g0396(.A1(new_n753_), .A2(G4092), .ZN(new_n762_));
  INV_X1    g0397(.A(new_n762_), .ZN(new_n763_));
  NOR3_X1   g0398(.A1(new_n760_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g0399(.A1(new_n757_), .A2(G129), .ZN(new_n765_));
  INV_X1    g0400(.A(KEYINPUT15), .ZN(new_n766_));
  NAND2_X1  g0401(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g0402(.A1(new_n757_), .A2(KEYINPUT15), .A3(G129), .ZN(new_n768_));
  AOI211_X1 g0403(.A(new_n759_), .B(new_n764_), .C1(new_n767_), .C2(new_n768_), .ZN(G838));
  INV_X1    g0404(.A(new_n587_), .ZN(new_n770_));
  NOR2_X1   g0405(.A1(new_n770_), .A2(new_n578_), .ZN(new_n771_));
  XOR2_X1   g0406(.A(new_n771_), .B(G4), .Z(new_n772_));
  OAI21_X1  g0407(.A(new_n756_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n773_));
  INV_X1    g0408(.A(G117), .ZN(new_n774_));
  AOI21_X1  g0409(.A(G4091), .B1(new_n774_), .B2(G4092), .ZN(new_n775_));
  AOI22_X1  g0410(.A1(new_n772_), .A2(new_n762_), .B1(new_n773_), .B2(new_n775_), .ZN(G861));
  OR2_X1    g0411(.A1(new_n661_), .A2(new_n747_), .ZN(new_n777_));
  NAND2_X1  g0412(.A1(new_n743_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g0413(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g0414(.A1(new_n673_), .A2(new_n736_), .ZN(new_n780_));
  NOR2_X1   g0415(.A1(new_n672_), .A2(new_n676_), .ZN(new_n781_));
  OAI211_X1 g0416(.A(new_n779_), .B(new_n780_), .C1(new_n686_), .C2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g0417(.A1(new_n682_), .A2(new_n676_), .ZN(new_n783_));
  XNOR2_X1  g0418(.A(new_n783_), .B(new_n686_), .ZN(new_n784_));
  OAI21_X1  g0419(.A(new_n782_), .B1(new_n779_), .B2(new_n784_), .ZN(G623));
  INV_X1    g0420(.A(G4087), .ZN(new_n786_));
  INV_X1    g0421(.A(G4088), .ZN(new_n787_));
  NOR2_X1   g0422(.A1(G861), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g0423(.A1(G822), .A2(G4088), .ZN(new_n789_));
  OAI21_X1  g0424(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g0425(.A1(G61), .A2(G4088), .ZN(new_n791_));
  INV_X1    g0426(.A(G11), .ZN(new_n792_));
  OAI21_X1  g0427(.A(new_n791_), .B1(new_n792_), .B2(G4088), .ZN(new_n793_));
  NAND2_X1  g0428(.A1(new_n793_), .A2(G4087), .ZN(new_n794_));
  NAND2_X1  g0429(.A1(new_n790_), .A2(new_n794_), .ZN(G722));
  NOR2_X1   g0430(.A1(new_n693_), .A2(new_n747_), .ZN(new_n796_));
  NAND2_X1  g0431(.A1(new_n648_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g0432(.A(new_n644_), .ZN(new_n798_));
  NOR2_X1   g0433(.A1(new_n798_), .A2(new_n640_), .ZN(new_n799_));
  AOI21_X1  g0434(.A(new_n660_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n800_));
  OAI211_X1 g0435(.A(new_n739_), .B(new_n799_), .C1(new_n800_), .C2(new_n629_), .ZN(new_n801_));
  NAND3_X1  g0436(.A1(new_n797_), .A2(new_n741_), .A3(new_n801_), .ZN(new_n802_));
  AOI22_X1  g0437(.A1(new_n802_), .A2(KEYINPUT16), .B1(new_n640_), .B2(new_n739_), .ZN(new_n803_));
  OAI21_X1  g0438(.A(new_n803_), .B1(KEYINPUT16), .B2(new_n802_), .ZN(new_n804_));
  XNOR2_X1  g0439(.A(new_n804_), .B(new_n696_), .ZN(new_n805_));
  NAND2_X1  g0440(.A1(new_n805_), .A2(new_n762_), .ZN(new_n806_));
  NAND2_X1  g0441(.A1(new_n465_), .A2(new_n756_), .ZN(new_n807_));
  OAI211_X1 g0442(.A(new_n807_), .B(new_n753_), .C1(G52), .C2(new_n756_), .ZN(new_n808_));
  NAND2_X1  g0443(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g0444(.A(new_n809_), .ZN(G832));
  OAI21_X1  g0445(.A(new_n644_), .B1(new_n760_), .B2(new_n629_), .ZN(new_n811_));
  NAND2_X1  g0446(.A1(new_n811_), .A2(new_n641_), .ZN(new_n812_));
  XNOR2_X1  g0447(.A(new_n812_), .B(new_n738_), .ZN(new_n813_));
  NAND2_X1  g0448(.A1(new_n813_), .A2(new_n762_), .ZN(new_n814_));
  NAND2_X1  g0449(.A1(G130), .A2(G4092), .ZN(new_n815_));
  OAI21_X1  g0450(.A(new_n815_), .B1(new_n467_), .B2(G4092), .ZN(new_n816_));
  NAND2_X1  g0451(.A1(new_n816_), .A2(new_n753_), .ZN(new_n817_));
  NAND2_X1  g0452(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g0453(.A(new_n818_), .ZN(G834));
  NOR2_X1   g0454(.A1(new_n457_), .A2(G4092), .ZN(new_n820_));
  NOR2_X1   g0455(.A1(new_n820_), .A2(KEYINPUT17), .ZN(new_n821_));
  AOI21_X1  g0456(.A(new_n821_), .B1(G119), .B2(G4092), .ZN(new_n822_));
  NAND2_X1  g0457(.A1(new_n820_), .A2(KEYINPUT17), .ZN(new_n823_));
  AOI21_X1  g0458(.A(G4091), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g0459(.A1(new_n632_), .A2(new_n660_), .A3(new_n625_), .ZN(new_n825_));
  AOI22_X1  g0460(.A1(new_n796_), .A2(new_n634_), .B1(new_n625_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g0461(.A(new_n826_), .B(new_n799_), .ZN(new_n827_));
  AOI21_X1  g0462(.A(new_n824_), .B1(new_n762_), .B2(new_n827_), .ZN(G836));
  INV_X1    g0463(.A(G4090), .ZN(new_n829_));
  INV_X1    g0464(.A(G4089), .ZN(new_n830_));
  NOR2_X1   g0465(.A1(G861), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g0466(.A1(G822), .A2(G4089), .ZN(new_n832_));
  OAI21_X1  g0467(.A(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g0468(.A1(G61), .A2(G4089), .ZN(new_n834_));
  OAI21_X1  g0469(.A(new_n834_), .B1(new_n792_), .B2(G4089), .ZN(new_n835_));
  NAND2_X1  g0470(.A1(new_n835_), .A2(G4090), .ZN(new_n836_));
  NAND2_X1  g0471(.A1(new_n833_), .A2(new_n836_), .ZN(G859));
  NAND2_X1  g0472(.A1(new_n589_), .A2(G4), .ZN(new_n838_));
  NAND2_X1  g0473(.A1(new_n838_), .A2(new_n727_), .ZN(new_n839_));
  INV_X1    g0474(.A(new_n586_), .ZN(new_n840_));
  NOR2_X1   g0475(.A1(new_n840_), .A2(new_n579_), .ZN(new_n841_));
  OAI21_X1  g0476(.A(new_n567_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g0477(.A(KEYINPUT18), .ZN(new_n843_));
  OAI221_X1 g0478(.A(new_n563_), .B1(new_n564_), .B2(new_n730_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g0479(.A(new_n844_), .B1(new_n843_), .B2(new_n842_), .ZN(new_n845_));
  XNOR2_X1  g0480(.A(new_n845_), .B(new_n574_), .ZN(new_n846_));
  OR2_X1    g0481(.A1(new_n846_), .A2(new_n763_), .ZN(new_n847_));
  NAND2_X1  g0482(.A1(new_n508_), .A2(new_n756_), .ZN(new_n848_));
  OAI211_X1 g0483(.A(new_n848_), .B(new_n753_), .C1(G122), .C2(new_n756_), .ZN(new_n849_));
  NAND2_X1  g0484(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g0485(.A(new_n850_), .ZN(G871));
  AOI21_X1  g0486(.A(new_n731_), .B1(new_n839_), .B2(new_n553_), .ZN(new_n852_));
  XNOR2_X1  g0487(.A(new_n852_), .B(new_n564_), .ZN(new_n853_));
  OR2_X1    g0488(.A1(new_n853_), .A2(new_n763_), .ZN(new_n854_));
  NAND2_X1  g0489(.A1(new_n495_), .A2(new_n756_), .ZN(new_n855_));
  OAI211_X1 g0490(.A(new_n855_), .B(new_n753_), .C1(G128), .C2(new_n756_), .ZN(new_n856_));
  NAND2_X1  g0491(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g0492(.A(new_n857_), .ZN(G873));
  OAI21_X1  g0493(.A(new_n753_), .B1(new_n756_), .B2(G127), .ZN(new_n859_));
  AOI21_X1  g0494(.A(new_n859_), .B1(new_n489_), .B2(new_n756_), .ZN(new_n860_));
  INV_X1    g0495(.A(new_n577_), .ZN(new_n861_));
  OAI211_X1 g0496(.A(new_n861_), .B(G374), .C1(new_n585_), .C2(KEYINPUT19), .ZN(new_n862_));
  AOI21_X1  g0497(.A(new_n862_), .B1(new_n840_), .B2(KEYINPUT19), .ZN(new_n863_));
  NOR2_X1   g0498(.A1(new_n839_), .A2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g0499(.A(new_n864_), .B(new_n556_), .ZN(new_n865_));
  AOI21_X1  g0500(.A(new_n860_), .B1(new_n865_), .B2(new_n762_), .ZN(G875));
  AOI21_X1  g0501(.A(new_n578_), .B1(G4), .B2(new_n587_), .ZN(new_n867_));
  XNOR2_X1  g0502(.A(new_n867_), .B(new_n586_), .ZN(new_n868_));
  OAI21_X1  g0503(.A(new_n756_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n869_));
  INV_X1    g0504(.A(G126), .ZN(new_n870_));
  AOI21_X1  g0505(.A(G4091), .B1(new_n870_), .B2(G4092), .ZN(new_n871_));
  AOI22_X1  g0506(.A1(new_n868_), .A2(new_n762_), .B1(new_n869_), .B2(new_n871_), .ZN(G877));
  NAND2_X1  g0507(.A1(new_n642_), .A2(new_n650_), .ZN(new_n873_));
  OAI21_X1  g0508(.A(new_n873_), .B1(G331), .B2(new_n642_), .ZN(new_n874_));
  XNOR2_X1  g0509(.A(new_n874_), .B(new_n639_), .ZN(new_n875_));
  MUX2_X1   g0510(.A(G369), .B(G372), .S(G332), .Z(new_n876_));
  XNOR2_X1  g0511(.A(new_n876_), .B(new_n660_), .ZN(new_n877_));
  XNOR2_X1  g0512(.A(new_n877_), .B(new_n631_), .ZN(new_n878_));
  XNOR2_X1  g0513(.A(new_n875_), .B(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g0514(.A(new_n879_), .B(new_n667_), .ZN(new_n880_));
  XNOR2_X1  g0515(.A(new_n685_), .B(new_n676_), .ZN(new_n881_));
  XNOR2_X1  g0516(.A(new_n881_), .B(new_n678_), .ZN(new_n882_));
  XNOR2_X1  g0517(.A(new_n882_), .B(KEYINPUT20), .ZN(new_n883_));
  XNOR2_X1  g0518(.A(new_n880_), .B(new_n883_), .ZN(G998));
  XNOR2_X1  g0519(.A(new_n577_), .B(new_n584_), .ZN(new_n885_));
  XNOR2_X1  g0520(.A(new_n885_), .B(new_n559_), .ZN(new_n886_));
  XNOR2_X1  g0521(.A(new_n886_), .B(new_n551_), .ZN(new_n887_));
  XOR2_X1   g0522(.A(new_n569_), .B(new_n593_), .Z(new_n888_));
  XNOR2_X1  g0523(.A(new_n888_), .B(new_n606_), .ZN(new_n889_));
  XNOR2_X1  g0524(.A(new_n887_), .B(new_n889_), .ZN(new_n890_));
  MUX2_X1   g0525(.A(G289), .B(G292), .S(G335), .Z(new_n891_));
  XNOR2_X1  g0526(.A(new_n600_), .B(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g0527(.A(new_n892_), .B(new_n613_), .ZN(new_n893_));
  XNOR2_X1  g0528(.A(new_n890_), .B(new_n893_), .ZN(G1000));
  NOR3_X1   g0529(.A1(new_n838_), .A2(new_n574_), .A3(new_n566_), .ZN(new_n895_));
  XOR2_X1   g0530(.A(new_n895_), .B(KEYINPUT21), .Z(new_n896_));
  INV_X1    g0531(.A(new_n734_), .ZN(new_n897_));
  NOR2_X1   g0532(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g0533(.A1(new_n619_), .A2(new_n596_), .ZN(new_n899_));
  NAND2_X1  g0534(.A1(new_n899_), .A2(new_n722_), .ZN(new_n900_));
  NAND2_X1  g0535(.A1(new_n900_), .A2(new_n609_), .ZN(new_n901_));
  NAND3_X1  g0536(.A1(new_n899_), .A2(new_n610_), .A3(new_n722_), .ZN(new_n902_));
  AOI21_X1  g0537(.A(new_n898_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g0538(.A(new_n898_), .B(KEYINPUT22), .ZN(new_n904_));
  NAND2_X1  g0539(.A1(new_n721_), .A2(new_n722_), .ZN(new_n905_));
  NAND2_X1  g0540(.A1(new_n905_), .A2(new_n609_), .ZN(new_n906_));
  NAND2_X1  g0541(.A1(new_n906_), .A2(new_n723_), .ZN(new_n907_));
  AOI21_X1  g0542(.A(new_n903_), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g0543(.A(KEYINPUT26), .ZN(new_n909_));
  AND2_X1   g0544(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g0545(.A(new_n724_), .B(new_n604_), .ZN(new_n911_));
  NAND2_X1  g0546(.A1(new_n904_), .A2(new_n911_), .ZN(new_n912_));
  XOR2_X1   g0547(.A(new_n604_), .B(KEYINPUT25), .Z(new_n913_));
  NAND2_X1  g0548(.A1(new_n902_), .A2(new_n607_), .ZN(new_n914_));
  XOR2_X1   g0549(.A(new_n913_), .B(new_n914_), .Z(new_n915_));
  OAI21_X1  g0550(.A(new_n912_), .B1(new_n898_), .B2(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g0551(.A(new_n898_), .B(new_n597_), .ZN(new_n917_));
  NOR3_X1   g0552(.A1(new_n865_), .A2(new_n772_), .A3(new_n868_), .ZN(new_n918_));
  NAND4_X1  g0553(.A1(new_n846_), .A2(new_n853_), .A3(new_n917_), .A4(new_n918_), .ZN(new_n919_));
  NOR3_X1   g0554(.A1(new_n910_), .A2(new_n916_), .A3(new_n919_), .ZN(new_n920_));
  OAI21_X1  g0555(.A(new_n920_), .B1(new_n909_), .B2(new_n908_), .ZN(new_n921_));
  OAI21_X1  g0556(.A(new_n595_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n922_));
  AND3_X1   g0557(.A1(new_n904_), .A2(new_n721_), .A3(new_n922_), .ZN(new_n923_));
  INV_X1    g0558(.A(KEYINPUT23), .ZN(new_n924_));
  OR2_X1    g0559(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g0560(.A1(new_n923_), .A2(new_n924_), .ZN(new_n926_));
  XNOR2_X1  g0561(.A(new_n619_), .B(new_n596_), .ZN(new_n927_));
  XNOR2_X1  g0562(.A(new_n927_), .B(KEYINPUT24), .ZN(new_n928_));
  OAI211_X1 g0563(.A(new_n925_), .B(new_n926_), .C1(new_n904_), .C2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g0564(.A1(new_n921_), .A2(new_n929_), .ZN(G575));
  MUX2_X1   g0565(.A(new_n672_), .B(new_n682_), .S(new_n778_), .Z(new_n931_));
  XNOR2_X1  g0566(.A(new_n931_), .B(new_n676_), .ZN(new_n932_));
  INV_X1    g0567(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g0568(.A1(new_n679_), .A2(new_n665_), .ZN(new_n934_));
  INV_X1    g0569(.A(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g0570(.A(new_n778_), .B(new_n935_), .ZN(new_n936_));
  INV_X1    g0571(.A(new_n668_), .ZN(new_n937_));
  NOR2_X1   g0572(.A1(new_n681_), .A2(new_n937_), .ZN(new_n938_));
  XOR2_X1   g0573(.A(new_n938_), .B(new_n665_), .Z(new_n939_));
  NAND2_X1  g0574(.A1(new_n779_), .A2(new_n939_), .ZN(new_n940_));
  NOR3_X1   g0575(.A1(new_n680_), .A2(new_n681_), .A3(new_n937_), .ZN(new_n941_));
  INV_X1    g0576(.A(new_n938_), .ZN(new_n942_));
  AOI21_X1  g0577(.A(new_n941_), .B1(new_n680_), .B2(new_n942_), .ZN(new_n943_));
  OAI21_X1  g0578(.A(new_n940_), .B1(new_n779_), .B2(new_n943_), .ZN(new_n944_));
  NAND4_X1  g0579(.A1(new_n933_), .A2(G623), .A3(new_n936_), .A4(new_n944_), .ZN(new_n945_));
  INV_X1    g0580(.A(KEYINPUT27), .ZN(new_n946_));
  AND2_X1   g0581(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g0582(.A1(new_n945_), .A2(new_n946_), .ZN(new_n948_));
  NAND3_X1  g0583(.A1(new_n634_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n949_));
  OR4_X1    g0584(.A1(new_n805_), .A2(new_n813_), .A3(new_n827_), .A4(new_n949_), .ZN(new_n950_));
  NOR3_X1   g0585(.A1(new_n947_), .A2(new_n948_), .A3(new_n950_), .ZN(G585));
  INV_X1    g0586(.A(G137), .ZN(new_n952_));
  INV_X1    g0587(.A(G1690), .ZN(new_n953_));
  INV_X1    g0588(.A(G1689), .ZN(new_n954_));
  NOR2_X1   g0589(.A1(G861), .A2(new_n954_), .ZN(new_n955_));
  NOR2_X1   g0590(.A1(G822), .A2(G1689), .ZN(new_n956_));
  OAI21_X1  g0591(.A(new_n953_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  MUX2_X1   g0592(.A(G182), .B(G185), .S(G1689), .Z(new_n958_));
  NAND2_X1  g0593(.A1(new_n958_), .A2(G1690), .ZN(new_n959_));
  AOI21_X1  g0594(.A(new_n952_), .B1(new_n957_), .B2(new_n959_), .ZN(G661));
  NOR2_X1   g0595(.A1(G822), .A2(G1694), .ZN(new_n961_));
  OR2_X1    g0596(.A1(new_n961_), .A2(KEYINPUT28), .ZN(new_n962_));
  AOI21_X1  g0597(.A(G1691), .B1(G182), .B2(G1694), .ZN(new_n963_));
  NAND2_X1  g0598(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  AOI21_X1  g0599(.A(new_n964_), .B1(KEYINPUT28), .B2(new_n961_), .ZN(new_n965_));
  INV_X1    g0600(.A(G1694), .ZN(new_n966_));
  NAND2_X1  g0601(.A1(G861), .A2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g0602(.A(new_n967_), .B1(G185), .B2(new_n966_), .ZN(new_n968_));
  AOI211_X1 g0603(.A(new_n952_), .B(new_n965_), .C1(G1691), .C2(new_n968_), .ZN(G693));
  NAND3_X1  g0604(.A1(new_n787_), .A2(G43), .A3(G4087), .ZN(new_n970_));
  NAND3_X1  g0605(.A1(G37), .A2(G4087), .A3(G4088), .ZN(new_n971_));
  XOR2_X1   g0606(.A(new_n971_), .B(KEYINPUT29), .Z(new_n972_));
  NOR2_X1   g0607(.A1(G832), .A2(G4088), .ZN(new_n973_));
  AOI21_X1  g0608(.A(new_n973_), .B1(new_n850_), .B2(G4088), .ZN(new_n974_));
  OAI211_X1 g0609(.A(new_n970_), .B(new_n972_), .C1(new_n974_), .C2(G4087), .ZN(new_n975_));
  XNOR2_X1  g0610(.A(new_n975_), .B(KEYINPUT30), .ZN(G747));
  NAND2_X1  g0611(.A1(new_n857_), .A2(new_n786_), .ZN(new_n977_));
  INV_X1    g0612(.A(KEYINPUT31), .ZN(new_n978_));
  NOR3_X1   g0613(.A1(new_n977_), .A2(new_n978_), .A3(new_n787_), .ZN(new_n979_));
  INV_X1    g0614(.A(G20), .ZN(new_n980_));
  OAI21_X1  g0615(.A(new_n977_), .B1(new_n980_), .B2(new_n786_), .ZN(new_n981_));
  AOI21_X1  g0616(.A(KEYINPUT31), .B1(new_n981_), .B2(G4088), .ZN(new_n982_));
  NOR2_X1   g0617(.A1(G834), .A2(G4087), .ZN(new_n983_));
  INV_X1    g0618(.A(G76), .ZN(new_n984_));
  NOR2_X1   g0619(.A1(new_n984_), .A2(new_n786_), .ZN(new_n985_));
  OAI21_X1  g0620(.A(new_n787_), .B1(new_n983_), .B2(new_n985_), .ZN(new_n986_));
  AOI21_X1  g0621(.A(new_n979_), .B1(new_n982_), .B2(new_n986_), .ZN(G752));
  NOR2_X1   g0622(.A1(G836), .A2(G4088), .ZN(new_n988_));
  NOR2_X1   g0623(.A1(G875), .A2(new_n787_), .ZN(new_n989_));
  OAI21_X1  g0624(.A(new_n786_), .B1(new_n988_), .B2(new_n989_), .ZN(new_n990_));
  NAND3_X1  g0625(.A1(new_n787_), .A2(G73), .A3(G4087), .ZN(new_n991_));
  NAND3_X1  g0626(.A1(G17), .A2(G4087), .A3(G4088), .ZN(new_n992_));
  XNOR2_X1  g0627(.A(new_n992_), .B(KEYINPUT32), .ZN(new_n993_));
  NAND3_X1  g0628(.A1(new_n990_), .A2(new_n991_), .A3(new_n993_), .ZN(G757));
  NOR2_X1   g0629(.A1(G838), .A2(G4088), .ZN(new_n995_));
  NOR2_X1   g0630(.A1(G877), .A2(new_n787_), .ZN(new_n996_));
  OAI21_X1  g0631(.A(new_n786_), .B1(new_n995_), .B2(new_n996_), .ZN(new_n997_));
  NAND2_X1  g0632(.A1(G70), .A2(G4088), .ZN(new_n998_));
  INV_X1    g0633(.A(G67), .ZN(new_n999_));
  OAI21_X1  g0634(.A(new_n998_), .B1(new_n999_), .B2(G4088), .ZN(new_n1000_));
  NAND2_X1  g0635(.A1(new_n1000_), .A2(G4087), .ZN(new_n1001_));
  NAND2_X1  g0636(.A1(new_n997_), .A2(new_n1001_), .ZN(G762));
  NOR2_X1   g0637(.A1(G871), .A2(new_n830_), .ZN(new_n1003_));
  NOR2_X1   g0638(.A1(G832), .A2(G4089), .ZN(new_n1004_));
  OAI21_X1  g0639(.A(new_n829_), .B1(new_n1003_), .B2(new_n1004_), .ZN(new_n1005_));
  INV_X1    g0640(.A(KEYINPUT33), .ZN(new_n1006_));
  MUX2_X1   g0641(.A(G43), .B(G37), .S(G4089), .Z(new_n1007_));
  AOI21_X1  g0642(.A(new_n1006_), .B1(new_n1007_), .B2(G4090), .ZN(new_n1008_));
  NOR2_X1   g0643(.A1(KEYINPUT33), .A2(G4090), .ZN(new_n1009_));
  AOI22_X1  g0644(.A1(new_n1005_), .A2(new_n1008_), .B1(new_n1003_), .B2(new_n1009_), .ZN(G787));
  NAND2_X1  g0645(.A1(G20), .A2(G4089), .ZN(new_n1011_));
  OAI21_X1  g0646(.A(new_n1011_), .B1(new_n984_), .B2(G4089), .ZN(new_n1012_));
  NAND2_X1  g0647(.A1(new_n1012_), .A2(G4090), .ZN(new_n1013_));
  NOR2_X1   g0648(.A1(G834), .A2(G4089), .ZN(new_n1014_));
  AOI21_X1  g0649(.A(new_n1014_), .B1(G4089), .B2(new_n857_), .ZN(new_n1015_));
  OAI21_X1  g0650(.A(new_n1013_), .B1(new_n1015_), .B2(G4090), .ZN(G792));
  NOR2_X1   g0651(.A1(G836), .A2(G4089), .ZN(new_n1017_));
  NOR2_X1   g0652(.A1(G875), .A2(new_n830_), .ZN(new_n1018_));
  OAI21_X1  g0653(.A(new_n829_), .B1(new_n1017_), .B2(new_n1018_), .ZN(new_n1019_));
  AND2_X1   g0654(.A1(G17), .A2(G4089), .ZN(new_n1020_));
  AOI21_X1  g0655(.A(new_n1020_), .B1(G73), .B2(new_n830_), .ZN(new_n1021_));
  OAI21_X1  g0656(.A(new_n1019_), .B1(new_n829_), .B2(new_n1021_), .ZN(G797));
  NOR2_X1   g0657(.A1(G838), .A2(G4089), .ZN(new_n1023_));
  NOR2_X1   g0658(.A1(G877), .A2(new_n830_), .ZN(new_n1024_));
  OAI21_X1  g0659(.A(new_n829_), .B1(new_n1023_), .B2(new_n1024_), .ZN(new_n1025_));
  NAND2_X1  g0660(.A1(G70), .A2(G4089), .ZN(new_n1026_));
  OAI21_X1  g0661(.A(new_n1026_), .B1(new_n999_), .B2(G4089), .ZN(new_n1027_));
  NAND2_X1  g0662(.A1(new_n1027_), .A2(G4090), .ZN(new_n1028_));
  NAND2_X1  g0663(.A1(new_n1025_), .A2(new_n1028_), .ZN(G802));
  NOR2_X1   g0664(.A1(G871), .A2(G1690), .ZN(new_n1030_));
  INV_X1    g0665(.A(G170), .ZN(new_n1031_));
  NOR2_X1   g0666(.A1(new_n1031_), .A2(new_n953_), .ZN(new_n1032_));
  OAI21_X1  g0667(.A(G1689), .B1(new_n1030_), .B2(new_n1032_), .ZN(new_n1033_));
  NOR2_X1   g0668(.A1(G832), .A2(G1690), .ZN(new_n1034_));
  INV_X1    g0669(.A(G200), .ZN(new_n1035_));
  NOR2_X1   g0670(.A1(new_n1035_), .A2(new_n953_), .ZN(new_n1036_));
  OAI21_X1  g0671(.A(new_n954_), .B1(new_n1034_), .B2(new_n1036_), .ZN(new_n1037_));
  AOI21_X1  g0672(.A(new_n952_), .B1(new_n1033_), .B2(new_n1037_), .ZN(G642));
  NOR2_X1   g0673(.A1(G838), .A2(G1690), .ZN(new_n1039_));
  INV_X1    g0674(.A(G188), .ZN(new_n1040_));
  NOR2_X1   g0675(.A1(new_n1040_), .A2(new_n953_), .ZN(new_n1041_));
  OAI21_X1  g0676(.A(new_n954_), .B1(new_n1039_), .B2(new_n1041_), .ZN(new_n1042_));
  NOR2_X1   g0677(.A1(G877), .A2(G1690), .ZN(new_n1043_));
  INV_X1    g0678(.A(G158), .ZN(new_n1044_));
  NOR2_X1   g0679(.A1(new_n1044_), .A2(new_n953_), .ZN(new_n1045_));
  OAI21_X1  g0680(.A(G1689), .B1(new_n1043_), .B2(new_n1045_), .ZN(new_n1046_));
  AOI21_X1  g0681(.A(new_n952_), .B1(new_n1042_), .B2(new_n1046_), .ZN(G664));
  NOR2_X1   g0682(.A1(G836), .A2(G1690), .ZN(new_n1048_));
  INV_X1    g0683(.A(G155), .ZN(new_n1049_));
  NOR2_X1   g0684(.A1(new_n1049_), .A2(new_n953_), .ZN(new_n1050_));
  OAI21_X1  g0685(.A(new_n954_), .B1(new_n1048_), .B2(new_n1050_), .ZN(new_n1051_));
  NOR2_X1   g0686(.A1(G875), .A2(G1690), .ZN(new_n1052_));
  INV_X1    g0687(.A(G152), .ZN(new_n1053_));
  NOR2_X1   g0688(.A1(new_n1053_), .A2(new_n953_), .ZN(new_n1054_));
  OAI21_X1  g0689(.A(G1689), .B1(new_n1052_), .B2(new_n1054_), .ZN(new_n1055_));
  AOI21_X1  g0690(.A(new_n952_), .B1(new_n1051_), .B2(new_n1055_), .ZN(G667));
  NAND3_X1  g0691(.A1(G146), .A2(G1689), .A3(G1690), .ZN(new_n1057_));
  INV_X1    g0692(.A(G149), .ZN(new_n1058_));
  NOR2_X1   g0693(.A1(new_n1058_), .A2(new_n953_), .ZN(new_n1059_));
  AOI21_X1  g0694(.A(new_n1059_), .B1(new_n818_), .B2(new_n953_), .ZN(new_n1060_));
  OAI21_X1  g0695(.A(new_n1057_), .B1(new_n1060_), .B2(G1689), .ZN(new_n1061_));
  OR2_X1    g0696(.A1(new_n1061_), .A2(KEYINPUT34), .ZN(new_n1062_));
  NOR2_X1   g0697(.A1(new_n954_), .A2(G1690), .ZN(new_n1063_));
  AOI22_X1  g0698(.A1(new_n1061_), .A2(KEYINPUT34), .B1(new_n857_), .B2(new_n1063_), .ZN(new_n1064_));
  AOI21_X1  g0699(.A(new_n952_), .B1(new_n1062_), .B2(new_n1064_), .ZN(G670));
  NOR2_X1   g0700(.A1(G871), .A2(G1694), .ZN(new_n1066_));
  NOR2_X1   g0701(.A1(new_n1031_), .A2(new_n966_), .ZN(new_n1067_));
  OAI21_X1  g0702(.A(G1691), .B1(new_n1066_), .B2(new_n1067_), .ZN(new_n1068_));
  INV_X1    g0703(.A(G1691), .ZN(new_n1069_));
  NOR2_X1   g0704(.A1(G832), .A2(G1694), .ZN(new_n1070_));
  NOR2_X1   g0705(.A1(new_n1035_), .A2(new_n966_), .ZN(new_n1071_));
  OAI21_X1  g0706(.A(new_n1069_), .B1(new_n1070_), .B2(new_n1071_), .ZN(new_n1072_));
  AOI21_X1  g0707(.A(new_n952_), .B1(new_n1068_), .B2(new_n1072_), .ZN(G676));
  NOR2_X1   g0708(.A1(G838), .A2(G1694), .ZN(new_n1074_));
  NOR2_X1   g0709(.A1(new_n1040_), .A2(new_n966_), .ZN(new_n1075_));
  OAI21_X1  g0710(.A(new_n1069_), .B1(new_n1074_), .B2(new_n1075_), .ZN(new_n1076_));
  NOR2_X1   g0711(.A1(G877), .A2(G1694), .ZN(new_n1077_));
  NOR2_X1   g0712(.A1(new_n1044_), .A2(new_n966_), .ZN(new_n1078_));
  OAI21_X1  g0713(.A(G1691), .B1(new_n1077_), .B2(new_n1078_), .ZN(new_n1079_));
  AOI21_X1  g0714(.A(new_n952_), .B1(new_n1076_), .B2(new_n1079_), .ZN(G696));
  NOR2_X1   g0715(.A1(G836), .A2(G1694), .ZN(new_n1081_));
  NOR2_X1   g0716(.A1(new_n1049_), .A2(new_n966_), .ZN(new_n1082_));
  OAI21_X1  g0717(.A(new_n1069_), .B1(new_n1081_), .B2(new_n1082_), .ZN(new_n1083_));
  NOR2_X1   g0718(.A1(G875), .A2(G1694), .ZN(new_n1084_));
  NOR2_X1   g0719(.A1(new_n1053_), .A2(new_n966_), .ZN(new_n1085_));
  OAI21_X1  g0720(.A(G1691), .B1(new_n1084_), .B2(new_n1085_), .ZN(new_n1086_));
  AOI21_X1  g0721(.A(new_n952_), .B1(new_n1083_), .B2(new_n1086_), .ZN(new_n1087_));
  XNOR2_X1  g0722(.A(new_n1087_), .B(KEYINPUT35), .ZN(G699));
  NOR2_X1   g0723(.A1(G834), .A2(G1694), .ZN(new_n1089_));
  NAND2_X1  g0724(.A1(new_n1089_), .A2(KEYINPUT37), .ZN(new_n1090_));
  INV_X1    g0725(.A(KEYINPUT37), .ZN(new_n1091_));
  OAI21_X1  g0726(.A(new_n1091_), .B1(new_n1058_), .B2(new_n966_), .ZN(new_n1092_));
  OAI211_X1 g0727(.A(new_n1090_), .B(new_n1069_), .C1(new_n1089_), .C2(new_n1092_), .ZN(new_n1093_));
  NAND3_X1  g0728(.A1(G146), .A2(G1691), .A3(G1694), .ZN(new_n1094_));
  XNOR2_X1  g0729(.A(new_n1094_), .B(KEYINPUT36), .ZN(new_n1095_));
  NOR2_X1   g0730(.A1(new_n1069_), .A2(G1694), .ZN(new_n1096_));
  AOI21_X1  g0731(.A(new_n1095_), .B1(new_n857_), .B2(new_n1096_), .ZN(new_n1097_));
  AOI21_X1  g0732(.A(new_n952_), .B1(new_n1093_), .B2(new_n1097_), .ZN(G702));
  NAND2_X1  g0733(.A1(G135), .A2(G4115), .ZN(new_n1099_));
  MUX2_X1   g0734(.A(new_n442_), .B(G123), .S(G3717), .Z(new_n1100_));
  OAI21_X1  g0735(.A(new_n1099_), .B1(new_n1100_), .B2(G3724), .ZN(new_n1101_));
  NAND2_X1  g0736(.A1(G623), .A2(G3717), .ZN(new_n1102_));
  XNOR2_X1  g0737(.A(new_n685_), .B(G132), .ZN(new_n1103_));
  OAI21_X1  g0738(.A(new_n1102_), .B1(G3717), .B2(new_n1103_), .ZN(new_n1104_));
  AOI21_X1  g0739(.A(new_n1101_), .B1(new_n1104_), .B2(G3724), .ZN(G818));
  XNOR2_X1  g0740(.A(G623), .B(new_n1103_), .ZN(G813));
  NAND2_X1  g0741(.A1(new_n442_), .A2(new_n753_), .ZN(new_n1107_));
  OAI21_X1  g0742(.A(new_n1107_), .B1(G623), .B2(new_n753_), .ZN(new_n1108_));
  AOI22_X1  g0743(.A1(new_n1108_), .A2(new_n756_), .B1(G123), .B2(new_n757_), .ZN(G824));
  NAND2_X1  g0744(.A1(G121), .A2(G4092), .ZN(new_n1110_));
  OAI21_X1  g0745(.A(new_n1110_), .B1(new_n445_), .B2(G4092), .ZN(new_n1111_));
  AOI22_X1  g0746(.A1(new_n932_), .A2(new_n762_), .B1(new_n753_), .B2(new_n1111_), .ZN(new_n1112_));
  XNOR2_X1  g0747(.A(new_n1112_), .B(KEYINPUT38), .ZN(G826));
  OR2_X1    g0748(.A1(new_n944_), .A2(new_n763_), .ZN(new_n1114_));
  OR2_X1    g0749(.A1(new_n432_), .A2(G4092), .ZN(new_n1115_));
  NAND2_X1  g0750(.A1(G116), .A2(G4092), .ZN(new_n1116_));
  XOR2_X1   g0751(.A(new_n1116_), .B(KEYINPUT39), .Z(new_n1117_));
  AOI21_X1  g0752(.A(G4091), .B1(new_n1115_), .B2(new_n1117_), .ZN(new_n1118_));
  XOR2_X1   g0753(.A(new_n1118_), .B(KEYINPUT40), .Z(new_n1119_));
  NAND2_X1  g0754(.A1(new_n1114_), .A2(new_n1119_), .ZN(new_n1120_));
  INV_X1    g0755(.A(new_n1120_), .ZN(G828));
  NAND2_X1  g0756(.A1(new_n757_), .A2(G112), .ZN(new_n1122_));
  MUX2_X1   g0757(.A(new_n439_), .B(new_n936_), .S(G4091), .Z(new_n1123_));
  OAI21_X1  g0758(.A(new_n1122_), .B1(new_n1123_), .B2(G4092), .ZN(new_n1124_));
  INV_X1    g0759(.A(new_n1124_), .ZN(G830));
  NAND4_X1  g0760(.A1(G245), .A2(G552), .A3(G559), .A4(G562), .ZN(new_n1126_));
  OR4_X1    g0761(.A1(G847), .A2(G1002), .A3(G1004), .A4(new_n1126_), .ZN(new_n1127_));
  NOR3_X1   g0762(.A1(G998), .A2(new_n1127_), .A3(G1000), .ZN(G854));
  NAND2_X1  g0763(.A1(new_n536_), .A2(new_n756_), .ZN(new_n1129_));
  NAND2_X1  g0764(.A1(G115), .A2(G4092), .ZN(new_n1130_));
  AOI21_X1  g0765(.A(G4091), .B1(new_n1129_), .B2(new_n1130_), .ZN(new_n1131_));
  AOI21_X1  g0766(.A(new_n1131_), .B1(new_n916_), .B2(new_n762_), .ZN(G863));
  NAND2_X1  g0767(.A1(new_n501_), .A2(new_n756_), .ZN(new_n1133_));
  OAI211_X1 g0768(.A(new_n1133_), .B(new_n753_), .C1(G114), .C2(new_n756_), .ZN(new_n1134_));
  OAI21_X1  g0769(.A(new_n1134_), .B1(new_n908_), .B2(new_n763_), .ZN(new_n1135_));
  XOR2_X1   g0770(.A(new_n1135_), .B(KEYINPUT41), .Z(G865));
  NAND2_X1  g0771(.A1(new_n929_), .A2(new_n762_), .ZN(new_n1137_));
  XOR2_X1   g0772(.A(new_n1137_), .B(KEYINPUT42), .Z(new_n1138_));
  OAI21_X1  g0773(.A(new_n753_), .B1(new_n756_), .B2(G53), .ZN(new_n1139_));
  AOI21_X1  g0774(.A(new_n1139_), .B1(new_n483_), .B2(new_n756_), .ZN(new_n1140_));
  NOR2_X1   g0775(.A1(new_n1138_), .A2(new_n1140_), .ZN(G867));
  OR2_X1    g0776(.A1(new_n917_), .A2(new_n763_), .ZN(new_n1142_));
  OR2_X1    g0777(.A1(new_n756_), .A2(G113), .ZN(new_n1143_));
  OAI211_X1 g0778(.A(new_n753_), .B(new_n1143_), .C1(new_n517_), .C2(G4092), .ZN(new_n1144_));
  NAND2_X1  g0779(.A1(new_n1142_), .A2(new_n1144_), .ZN(new_n1145_));
  INV_X1    g0780(.A(new_n1145_), .ZN(G869));
  NAND2_X1  g0781(.A1(G106), .A2(G4089), .ZN(new_n1147_));
  INV_X1    g0782(.A(G109), .ZN(new_n1148_));
  OAI21_X1  g0783(.A(new_n1147_), .B1(new_n1148_), .B2(G4089), .ZN(new_n1149_));
  NAND2_X1  g0784(.A1(new_n1149_), .A2(G4090), .ZN(new_n1150_));
  NOR2_X1   g0785(.A1(G824), .A2(G4089), .ZN(new_n1151_));
  XOR2_X1   g0786(.A(G863), .B(KEYINPUT43), .Z(new_n1152_));
  AOI21_X1  g0787(.A(new_n1151_), .B1(new_n1152_), .B2(G4089), .ZN(new_n1153_));
  OAI21_X1  g0788(.A(new_n1150_), .B1(new_n1153_), .B2(G4090), .ZN(G712));
  NAND2_X1  g0789(.A1(G106), .A2(G4088), .ZN(new_n1155_));
  OAI21_X1  g0790(.A(new_n1155_), .B1(new_n1148_), .B2(G4088), .ZN(new_n1156_));
  NAND2_X1  g0791(.A1(new_n1156_), .A2(G4087), .ZN(new_n1157_));
  NOR2_X1   g0792(.A1(G824), .A2(G4088), .ZN(new_n1158_));
  AOI21_X1  g0793(.A(new_n1158_), .B1(new_n1152_), .B2(G4088), .ZN(new_n1159_));
  OAI21_X1  g0794(.A(new_n1157_), .B1(new_n1159_), .B2(G4087), .ZN(G727));
  NOR2_X1   g0795(.A1(G826), .A2(G4088), .ZN(new_n1161_));
  NOR2_X1   g0796(.A1(G865), .A2(new_n787_), .ZN(new_n1162_));
  OAI21_X1  g0797(.A(new_n786_), .B1(new_n1161_), .B2(new_n1162_), .ZN(new_n1163_));
  NAND2_X1  g0798(.A1(G49), .A2(G4088), .ZN(new_n1164_));
  INV_X1    g0799(.A(G46), .ZN(new_n1165_));
  OAI21_X1  g0800(.A(new_n1164_), .B1(new_n1165_), .B2(G4088), .ZN(new_n1166_));
  NAND2_X1  g0801(.A1(new_n1166_), .A2(G4087), .ZN(new_n1167_));
  NAND2_X1  g0802(.A1(new_n1163_), .A2(new_n1167_), .ZN(G732));
  NAND2_X1  g0803(.A1(G103), .A2(G4088), .ZN(new_n1169_));
  INV_X1    g0804(.A(G100), .ZN(new_n1170_));
  OAI21_X1  g0805(.A(new_n1169_), .B1(new_n1170_), .B2(G4088), .ZN(new_n1171_));
  NAND2_X1  g0806(.A1(new_n1171_), .A2(G4087), .ZN(new_n1172_));
  MUX2_X1   g0807(.A(G828), .B(G867), .S(G4088), .Z(new_n1173_));
  OAI21_X1  g0808(.A(new_n1172_), .B1(new_n1173_), .B2(G4087), .ZN(G737));
  NAND2_X1  g0809(.A1(G40), .A2(G4088), .ZN(new_n1175_));
  INV_X1    g0810(.A(G91), .ZN(new_n1176_));
  OAI21_X1  g0811(.A(new_n1175_), .B1(new_n1176_), .B2(G4088), .ZN(new_n1177_));
  NAND2_X1  g0812(.A1(new_n1177_), .A2(G4087), .ZN(new_n1178_));
  MUX2_X1   g0813(.A(G830), .B(G869), .S(G4088), .Z(new_n1179_));
  OAI21_X1  g0814(.A(new_n1178_), .B1(new_n1179_), .B2(G4087), .ZN(G742));
  NOR2_X1   g0815(.A1(G826), .A2(G4089), .ZN(new_n1181_));
  NOR2_X1   g0816(.A1(G865), .A2(new_n830_), .ZN(new_n1182_));
  OAI21_X1  g0817(.A(new_n829_), .B1(new_n1181_), .B2(new_n1182_), .ZN(new_n1183_));
  NAND2_X1  g0818(.A1(G49), .A2(G4089), .ZN(new_n1184_));
  OAI21_X1  g0819(.A(new_n1184_), .B1(new_n1165_), .B2(G4089), .ZN(new_n1185_));
  NAND2_X1  g0820(.A1(new_n1185_), .A2(G4090), .ZN(new_n1186_));
  NAND2_X1  g0821(.A1(new_n1183_), .A2(new_n1186_), .ZN(G772));
  NAND2_X1  g0822(.A1(G103), .A2(G4089), .ZN(new_n1188_));
  OAI21_X1  g0823(.A(new_n1188_), .B1(new_n1170_), .B2(G4089), .ZN(new_n1189_));
  NAND2_X1  g0824(.A1(new_n1189_), .A2(G4090), .ZN(new_n1190_));
  MUX2_X1   g0825(.A(G828), .B(G867), .S(G4089), .Z(new_n1191_));
  OAI21_X1  g0826(.A(new_n1190_), .B1(new_n1191_), .B2(G4090), .ZN(G777));
  NAND2_X1  g0827(.A1(G40), .A2(G4089), .ZN(new_n1193_));
  OAI21_X1  g0828(.A(new_n1193_), .B1(new_n1176_), .B2(G4089), .ZN(new_n1194_));
  NAND2_X1  g0829(.A1(new_n1194_), .A2(G4090), .ZN(new_n1195_));
  MUX2_X1   g0830(.A(G830), .B(G869), .S(G4089), .Z(new_n1196_));
  OAI21_X1  g0831(.A(new_n1195_), .B1(new_n1196_), .B2(G4090), .ZN(G782));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1198_));
  INV_X1    g0833(.A(G203), .ZN(new_n1199_));
  OAI21_X1  g0834(.A(new_n1198_), .B1(new_n1199_), .B2(new_n953_), .ZN(new_n1200_));
  NAND3_X1  g0835(.A1(KEYINPUT45), .A2(G203), .A3(G1690), .ZN(new_n1201_));
  NAND3_X1  g0836(.A1(new_n1200_), .A2(new_n954_), .A3(new_n1201_), .ZN(new_n1202_));
  NAND3_X1  g0837(.A1(G173), .A2(G1689), .A3(G1690), .ZN(new_n1203_));
  NAND2_X1  g0838(.A1(new_n1203_), .A2(KEYINPUT44), .ZN(new_n1204_));
  OR2_X1    g0839(.A1(new_n1203_), .A2(KEYINPUT44), .ZN(new_n1205_));
  NAND3_X1  g0840(.A1(new_n1202_), .A2(new_n1204_), .A3(new_n1205_), .ZN(new_n1206_));
  AOI21_X1  g0841(.A(new_n1206_), .B1(new_n1145_), .B2(new_n1063_), .ZN(new_n1207_));
  NAND3_X1  g0842(.A1(new_n1124_), .A2(new_n954_), .A3(new_n953_), .ZN(new_n1208_));
  AOI21_X1  g0843(.A(new_n952_), .B1(new_n1207_), .B2(new_n1208_), .ZN(G645));
  NAND2_X1  g0844(.A1(new_n1120_), .A2(new_n954_), .ZN(new_n1210_));
  OAI21_X1  g0845(.A(new_n1210_), .B1(G867), .B2(new_n954_), .ZN(new_n1211_));
  NAND2_X1  g0846(.A1(new_n1211_), .A2(new_n953_), .ZN(new_n1212_));
  NAND2_X1  g0847(.A1(G167), .A2(G1689), .ZN(new_n1213_));
  INV_X1    g0848(.A(G197), .ZN(new_n1214_));
  OAI21_X1  g0849(.A(new_n1213_), .B1(new_n1214_), .B2(G1689), .ZN(new_n1215_));
  NAND2_X1  g0850(.A1(new_n1215_), .A2(G1690), .ZN(new_n1216_));
  AOI21_X1  g0851(.A(new_n952_), .B1(new_n1212_), .B2(new_n1216_), .ZN(G648));
  NOR2_X1   g0852(.A1(G826), .A2(G1690), .ZN(new_n1218_));
  INV_X1    g0853(.A(G194), .ZN(new_n1219_));
  NOR2_X1   g0854(.A1(new_n1219_), .A2(new_n953_), .ZN(new_n1220_));
  OAI21_X1  g0855(.A(new_n954_), .B1(new_n1218_), .B2(new_n1220_), .ZN(new_n1221_));
  NAND2_X1  g0856(.A1(G164), .A2(G1690), .ZN(new_n1222_));
  OAI21_X1  g0857(.A(new_n1222_), .B1(G865), .B2(G1690), .ZN(new_n1223_));
  NAND2_X1  g0858(.A1(new_n1223_), .A2(G1689), .ZN(new_n1224_));
  AOI21_X1  g0859(.A(new_n952_), .B1(new_n1221_), .B2(new_n1224_), .ZN(G651));
  AND2_X1   g0860(.A1(new_n1152_), .A2(new_n953_), .ZN(new_n1226_));
  INV_X1    g0861(.A(G161), .ZN(new_n1227_));
  NOR2_X1   g0862(.A1(new_n1227_), .A2(new_n953_), .ZN(new_n1228_));
  OAI21_X1  g0863(.A(G1689), .B1(new_n1226_), .B2(new_n1228_), .ZN(new_n1229_));
  NAND2_X1  g0864(.A1(G191), .A2(G1690), .ZN(new_n1230_));
  OAI21_X1  g0865(.A(new_n1230_), .B1(G824), .B2(G1690), .ZN(new_n1231_));
  NAND2_X1  g0866(.A1(new_n1231_), .A2(new_n954_), .ZN(new_n1232_));
  AOI21_X1  g0867(.A(new_n952_), .B1(new_n1229_), .B2(new_n1232_), .ZN(G654));
  NOR2_X1   g0868(.A1(G869), .A2(G1694), .ZN(new_n1234_));
  AND2_X1   g0869(.A1(G173), .A2(G1694), .ZN(new_n1235_));
  OAI21_X1  g0870(.A(G1691), .B1(new_n1234_), .B2(new_n1235_), .ZN(new_n1236_));
  NOR2_X1   g0871(.A1(G830), .A2(G1694), .ZN(new_n1237_));
  NOR2_X1   g0872(.A1(new_n1199_), .A2(new_n966_), .ZN(new_n1238_));
  OAI21_X1  g0873(.A(new_n1069_), .B1(new_n1237_), .B2(new_n1238_), .ZN(new_n1239_));
  AOI21_X1  g0874(.A(new_n952_), .B1(new_n1236_), .B2(new_n1239_), .ZN(G679));
  NAND2_X1  g0875(.A1(new_n1120_), .A2(new_n1069_), .ZN(new_n1241_));
  OAI21_X1  g0876(.A(new_n1241_), .B1(G867), .B2(new_n1069_), .ZN(new_n1242_));
  NAND2_X1  g0877(.A1(new_n1242_), .A2(new_n966_), .ZN(new_n1243_));
  NAND2_X1  g0878(.A1(G167), .A2(G1691), .ZN(new_n1244_));
  OAI21_X1  g0879(.A(new_n1244_), .B1(new_n1214_), .B2(G1691), .ZN(new_n1245_));
  NAND2_X1  g0880(.A1(new_n1245_), .A2(G1694), .ZN(new_n1246_));
  AOI21_X1  g0881(.A(new_n952_), .B1(new_n1243_), .B2(new_n1246_), .ZN(G682));
  NOR2_X1   g0882(.A1(G826), .A2(G1694), .ZN(new_n1248_));
  NOR2_X1   g0883(.A1(new_n1219_), .A2(new_n966_), .ZN(new_n1249_));
  OAI21_X1  g0884(.A(new_n1069_), .B1(new_n1248_), .B2(new_n1249_), .ZN(new_n1250_));
  NAND2_X1  g0885(.A1(G164), .A2(G1694), .ZN(new_n1251_));
  OAI21_X1  g0886(.A(new_n1251_), .B1(G865), .B2(G1694), .ZN(new_n1252_));
  NAND2_X1  g0887(.A1(new_n1252_), .A2(G1691), .ZN(new_n1253_));
  AOI21_X1  g0888(.A(new_n952_), .B1(new_n1250_), .B2(new_n1253_), .ZN(G685));
  AND2_X1   g0889(.A1(new_n1152_), .A2(new_n966_), .ZN(new_n1255_));
  NOR2_X1   g0890(.A1(new_n1227_), .A2(new_n966_), .ZN(new_n1256_));
  OAI21_X1  g0891(.A(G1691), .B1(new_n1255_), .B2(new_n1256_), .ZN(new_n1257_));
  NAND2_X1  g0892(.A1(G191), .A2(G1694), .ZN(new_n1258_));
  OAI21_X1  g0893(.A(new_n1258_), .B1(G824), .B2(G1694), .ZN(new_n1259_));
  NAND2_X1  g0894(.A1(new_n1259_), .A2(new_n1069_), .ZN(new_n1260_));
  AOI21_X1  g0895(.A(new_n952_), .B1(new_n1257_), .B2(new_n1260_), .ZN(G688));
  OAI21_X1  g0896(.A(G4092), .B1(G120), .B2(G4091), .ZN(new_n1262_));
  NOR3_X1   g0897(.A1(new_n626_), .A2(new_n629_), .A3(new_n622_), .ZN(new_n1263_));
  AOI21_X1  g0898(.A(KEYINPUT10), .B1(new_n632_), .B2(new_n625_), .ZN(new_n1264_));
  OAI21_X1  g0899(.A(new_n659_), .B1(new_n1263_), .B2(new_n1264_), .ZN(new_n1265_));
  AOI21_X1  g0900(.A(KEYINPUT47), .B1(new_n1265_), .B2(new_n632_), .ZN(new_n1266_));
  INV_X1    g0901(.A(KEYINPUT47), .ZN(new_n1267_));
  NOR3_X1   g0902(.A1(new_n800_), .A2(new_n1267_), .A3(new_n629_), .ZN(new_n1268_));
  INV_X1    g0903(.A(KEYINPUT11), .ZN(new_n1269_));
  NAND2_X1  g0904(.A1(new_n659_), .A2(new_n1269_), .ZN(new_n1270_));
  AOI21_X1  g0905(.A(new_n629_), .B1(new_n1270_), .B2(new_n690_), .ZN(new_n1271_));
  OAI21_X1  g0906(.A(new_n641_), .B1(new_n1271_), .B2(new_n626_), .ZN(new_n1272_));
  AOI21_X1  g0907(.A(new_n693_), .B1(new_n1272_), .B2(new_n644_), .ZN(new_n1273_));
  NAND3_X1  g0908(.A1(new_n825_), .A2(new_n644_), .A3(new_n625_), .ZN(new_n1274_));
  AOI21_X1  g0909(.A(new_n660_), .B1(new_n1274_), .B2(new_n641_), .ZN(new_n1275_));
  OAI22_X1  g0910(.A1(new_n1266_), .A2(new_n1268_), .B1(new_n1273_), .B2(new_n1275_), .ZN(new_n1276_));
  OAI21_X1  g0911(.A(new_n632_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n1277_));
  AOI21_X1  g0912(.A(new_n640_), .B1(new_n1277_), .B2(new_n625_), .ZN(new_n1278_));
  OAI21_X1  g0913(.A(new_n694_), .B1(new_n1278_), .B2(new_n798_), .ZN(new_n1279_));
  OAI21_X1  g0914(.A(new_n1267_), .B1(new_n800_), .B2(new_n629_), .ZN(new_n1280_));
  NAND3_X1  g0915(.A1(new_n1265_), .A2(KEYINPUT47), .A3(new_n632_), .ZN(new_n1281_));
  NAND2_X1  g0916(.A1(new_n1274_), .A2(new_n641_), .ZN(new_n1282_));
  NAND2_X1  g0917(.A1(new_n1282_), .A2(new_n659_), .ZN(new_n1283_));
  NAND4_X1  g0918(.A1(new_n1279_), .A2(new_n1280_), .A3(new_n1281_), .A4(new_n1283_), .ZN(new_n1284_));
  NAND3_X1  g0919(.A1(new_n1276_), .A2(KEYINPUT48), .A3(new_n1284_), .ZN(new_n1285_));
  NAND3_X1  g0920(.A1(new_n643_), .A2(new_n640_), .A3(new_n646_), .ZN(new_n1286_));
  AOI21_X1  g0921(.A(new_n629_), .B1(new_n634_), .B2(new_n659_), .ZN(new_n1287_));
  OAI211_X1 g0922(.A(new_n741_), .B(new_n1286_), .C1(new_n1287_), .C2(new_n647_), .ZN(new_n1288_));
  INV_X1    g0923(.A(KEYINPUT46), .ZN(new_n1289_));
  NAND2_X1  g0924(.A1(new_n1288_), .A2(new_n1289_), .ZN(new_n1290_));
  NAND4_X1  g0925(.A1(new_n801_), .A2(KEYINPUT46), .A3(new_n741_), .A4(new_n1286_), .ZN(new_n1291_));
  NOR2_X1   g0926(.A1(new_n1266_), .A2(new_n1268_), .ZN(new_n1292_));
  INV_X1    g0927(.A(KEYINPUT48), .ZN(new_n1293_));
  NOR2_X1   g0928(.A1(new_n1273_), .A2(new_n1275_), .ZN(new_n1294_));
  NAND3_X1  g0929(.A1(new_n1292_), .A2(new_n1293_), .A3(new_n1294_), .ZN(new_n1295_));
  NAND4_X1  g0930(.A1(new_n1285_), .A2(new_n1290_), .A3(new_n1291_), .A4(new_n1295_), .ZN(new_n1296_));
  NAND2_X1  g0931(.A1(new_n1290_), .A2(new_n1291_), .ZN(new_n1297_));
  NAND2_X1  g0932(.A1(new_n1277_), .A2(new_n625_), .ZN(new_n1298_));
  NAND3_X1  g0933(.A1(new_n1272_), .A2(new_n644_), .A3(new_n693_), .ZN(new_n1299_));
  NAND3_X1  g0934(.A1(new_n1274_), .A2(new_n641_), .A3(new_n660_), .ZN(new_n1300_));
  AOI21_X1  g0935(.A(new_n1298_), .B1(new_n1299_), .B2(new_n1300_), .ZN(new_n1301_));
  AOI21_X1  g0936(.A(new_n1301_), .B1(new_n1292_), .B2(new_n1294_), .ZN(new_n1302_));
  AOI21_X1  g0937(.A(new_n660_), .B1(new_n1297_), .B2(new_n1302_), .ZN(new_n1303_));
  NAND2_X1  g0938(.A1(new_n1296_), .A2(new_n1303_), .ZN(new_n1304_));
  INV_X1    g0939(.A(KEYINPUT49), .ZN(new_n1305_));
  NAND2_X1  g0940(.A1(new_n1304_), .A2(new_n1305_), .ZN(new_n1306_));
  NAND3_X1  g0941(.A1(new_n1296_), .A2(new_n1303_), .A3(KEYINPUT49), .ZN(new_n1307_));
  NAND2_X1  g0942(.A1(new_n1306_), .A2(new_n1307_), .ZN(new_n1308_));
  AOI22_X1  g0943(.A1(new_n1285_), .A2(new_n1295_), .B1(new_n1290_), .B2(new_n1291_), .ZN(new_n1309_));
  NOR2_X1   g0944(.A1(new_n1297_), .A2(new_n1302_), .ZN(new_n1310_));
  OAI21_X1  g0945(.A(new_n694_), .B1(new_n1309_), .B2(new_n1310_), .ZN(new_n1311_));
  AOI21_X1  g0946(.A(new_n635_), .B1(new_n1308_), .B2(new_n1311_), .ZN(new_n1312_));
  NAND2_X1  g0947(.A1(new_n1285_), .A2(new_n1295_), .ZN(new_n1313_));
  NAND2_X1  g0948(.A1(new_n1313_), .A2(new_n1297_), .ZN(new_n1314_));
  OR2_X1    g0949(.A1(new_n1297_), .A2(new_n1302_), .ZN(new_n1315_));
  AOI21_X1  g0950(.A(new_n693_), .B1(new_n1314_), .B2(new_n1315_), .ZN(new_n1316_));
  NOR3_X1   g0951(.A1(new_n1309_), .A2(new_n1310_), .A3(new_n694_), .ZN(new_n1317_));
  NOR3_X1   g0952(.A1(new_n1316_), .A2(new_n1317_), .A3(new_n634_), .ZN(new_n1318_));
  NOR3_X1   g0953(.A1(new_n1312_), .A2(new_n656_), .A3(new_n1318_), .ZN(new_n1319_));
  AND3_X1   g0954(.A1(new_n1296_), .A2(new_n1303_), .A3(KEYINPUT49), .ZN(new_n1320_));
  AOI21_X1  g0955(.A(KEYINPUT49), .B1(new_n1296_), .B2(new_n1303_), .ZN(new_n1321_));
  OAI21_X1  g0956(.A(new_n1311_), .B1(new_n1320_), .B2(new_n1321_), .ZN(new_n1322_));
  NAND2_X1  g0957(.A1(new_n1322_), .A2(new_n634_), .ZN(new_n1323_));
  OR3_X1    g0958(.A1(new_n1316_), .A2(new_n1317_), .A3(new_n634_), .ZN(new_n1324_));
  AOI21_X1  g0959(.A(new_n696_), .B1(new_n1323_), .B2(new_n1324_), .ZN(new_n1325_));
  OAI21_X1  g0960(.A(new_n799_), .B1(new_n1319_), .B2(new_n1325_), .ZN(new_n1326_));
  OAI21_X1  g0961(.A(new_n656_), .B1(new_n1312_), .B2(new_n1318_), .ZN(new_n1327_));
  OAI211_X1 g0962(.A(new_n635_), .B(new_n1311_), .C1(new_n1320_), .C2(new_n1321_), .ZN(new_n1328_));
  OAI21_X1  g0963(.A(new_n634_), .B1(new_n1316_), .B2(new_n1317_), .ZN(new_n1329_));
  NAND3_X1  g0964(.A1(new_n1328_), .A2(new_n1329_), .A3(new_n696_), .ZN(new_n1330_));
  INV_X1    g0965(.A(KEYINPUT50), .ZN(new_n1331_));
  NAND2_X1  g0966(.A1(new_n1330_), .A2(new_n1331_), .ZN(new_n1332_));
  INV_X1    g0967(.A(new_n799_), .ZN(new_n1333_));
  NAND4_X1  g0968(.A1(new_n1328_), .A2(new_n1329_), .A3(KEYINPUT50), .A4(new_n696_), .ZN(new_n1334_));
  NAND4_X1  g0969(.A1(new_n1327_), .A2(new_n1332_), .A3(new_n1333_), .A4(new_n1334_), .ZN(new_n1335_));
  NAND3_X1  g0970(.A1(new_n1326_), .A2(new_n1335_), .A3(new_n738_), .ZN(new_n1336_));
  OAI21_X1  g0971(.A(new_n1333_), .B1(new_n1319_), .B2(new_n1325_), .ZN(new_n1337_));
  NAND4_X1  g0972(.A1(new_n1327_), .A2(new_n1332_), .A3(new_n799_), .A4(new_n1334_), .ZN(new_n1338_));
  NAND3_X1  g0973(.A1(new_n1337_), .A2(new_n1338_), .A3(new_n739_), .ZN(new_n1339_));
  INV_X1    g0974(.A(G2174), .ZN(new_n1340_));
  NAND3_X1  g0975(.A1(new_n1336_), .A2(new_n1339_), .A3(new_n1340_), .ZN(new_n1341_));
  NAND3_X1  g0976(.A1(new_n1298_), .A2(new_n640_), .A3(new_n825_), .ZN(new_n1342_));
  XOR2_X1   g0977(.A(new_n1342_), .B(KEYINPUT51), .Z(new_n1343_));
  NAND2_X1  g0978(.A1(new_n1292_), .A2(new_n825_), .ZN(new_n1344_));
  NAND2_X1  g0979(.A1(new_n1298_), .A2(new_n825_), .ZN(new_n1345_));
  AOI21_X1  g0980(.A(new_n640_), .B1(new_n1345_), .B2(new_n644_), .ZN(new_n1346_));
  AOI21_X1  g0981(.A(new_n1343_), .B1(new_n1344_), .B2(new_n1346_), .ZN(new_n1347_));
  NAND4_X1  g0982(.A1(new_n695_), .A2(new_n741_), .A3(new_n801_), .A4(new_n1286_), .ZN(new_n1348_));
  NOR2_X1   g0983(.A1(new_n1347_), .A2(new_n1348_), .ZN(new_n1349_));
  NAND2_X1  g0984(.A1(new_n1347_), .A2(new_n1348_), .ZN(new_n1350_));
  INV_X1    g0985(.A(KEYINPUT52), .ZN(new_n1351_));
  NAND2_X1  g0986(.A1(new_n1350_), .A2(new_n1351_), .ZN(new_n1352_));
  NAND3_X1  g0987(.A1(new_n1347_), .A2(KEYINPUT52), .A3(new_n1348_), .ZN(new_n1353_));
  AOI21_X1  g0988(.A(new_n1349_), .B1(new_n1352_), .B2(new_n1353_), .ZN(new_n1354_));
  OAI21_X1  g0989(.A(new_n634_), .B1(new_n1354_), .B2(new_n1269_), .ZN(new_n1355_));
  INV_X1    g0990(.A(new_n1355_), .ZN(new_n1356_));
  NOR2_X1   g0991(.A1(new_n1354_), .A2(new_n634_), .ZN(new_n1357_));
  OAI21_X1  g0992(.A(new_n694_), .B1(new_n1356_), .B2(new_n1357_), .ZN(new_n1358_));
  OAI211_X1 g0993(.A(new_n1355_), .B(new_n693_), .C1(new_n634_), .C2(new_n1354_), .ZN(new_n1359_));
  NAND2_X1  g0994(.A1(new_n1358_), .A2(new_n1359_), .ZN(new_n1360_));
  XOR2_X1   g0995(.A(new_n799_), .B(new_n656_), .Z(new_n1361_));
  XNOR2_X1  g0996(.A(new_n1361_), .B(new_n738_), .ZN(new_n1362_));
  INV_X1    g0997(.A(new_n1362_), .ZN(new_n1363_));
  NAND2_X1  g0998(.A1(new_n1360_), .A2(new_n1363_), .ZN(new_n1364_));
  NAND3_X1  g0999(.A1(new_n1358_), .A2(new_n1362_), .A3(new_n1359_), .ZN(new_n1365_));
  NAND3_X1  g1000(.A1(new_n1364_), .A2(G2174), .A3(new_n1365_), .ZN(new_n1366_));
  NAND2_X1  g1001(.A1(new_n1341_), .A2(new_n1366_), .ZN(new_n1367_));
  AOI21_X1  g1002(.A(new_n942_), .B1(new_n781_), .B2(new_n935_), .ZN(new_n1368_));
  NAND2_X1  g1003(.A1(new_n781_), .A2(new_n669_), .ZN(new_n1369_));
  XOR2_X1   g1004(.A(new_n1369_), .B(KEYINPUT54), .Z(new_n1370_));
  OAI21_X1  g1005(.A(new_n680_), .B1(new_n677_), .B2(new_n937_), .ZN(new_n1371_));
  NAND3_X1  g1006(.A1(new_n681_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n1372_));
  AOI21_X1  g1007(.A(new_n935_), .B1(new_n1371_), .B2(new_n1372_), .ZN(new_n1373_));
  AND2_X1   g1008(.A1(new_n935_), .A2(new_n1372_), .ZN(new_n1374_));
  NOR2_X1   g1009(.A1(new_n1373_), .A2(new_n1374_), .ZN(new_n1375_));
  OAI22_X1  g1010(.A1(new_n1375_), .A2(new_n938_), .B1(new_n676_), .B2(new_n672_), .ZN(new_n1376_));
  AND2_X1   g1011(.A1(new_n1370_), .A2(new_n1376_), .ZN(new_n1377_));
  OAI21_X1  g1012(.A(new_n1368_), .B1(new_n1377_), .B2(new_n935_), .ZN(new_n1378_));
  INV_X1    g1013(.A(KEYINPUT55), .ZN(new_n1379_));
  XNOR2_X1  g1014(.A(new_n1378_), .B(new_n1379_), .ZN(new_n1380_));
  NOR2_X1   g1015(.A1(new_n1373_), .A2(new_n938_), .ZN(new_n1381_));
  OAI21_X1  g1016(.A(new_n1381_), .B1(new_n1377_), .B2(new_n934_), .ZN(new_n1382_));
  NAND3_X1  g1017(.A1(new_n1380_), .A2(new_n677_), .A3(new_n1382_), .ZN(new_n1383_));
  INV_X1    g1018(.A(new_n1383_), .ZN(new_n1384_));
  AOI21_X1  g1019(.A(new_n677_), .B1(new_n1380_), .B2(new_n1382_), .ZN(new_n1385_));
  OAI21_X1  g1020(.A(new_n686_), .B1(new_n1384_), .B2(new_n1385_), .ZN(new_n1386_));
  INV_X1    g1021(.A(new_n1385_), .ZN(new_n1387_));
  NAND3_X1  g1022(.A1(new_n1387_), .A2(new_n685_), .A3(new_n1383_), .ZN(new_n1388_));
  OAI21_X1  g1023(.A(new_n743_), .B1(new_n1340_), .B2(new_n698_), .ZN(new_n1389_));
  INV_X1    g1024(.A(new_n1389_), .ZN(new_n1390_));
  NAND3_X1  g1025(.A1(new_n1386_), .A2(new_n1388_), .A3(new_n1390_), .ZN(new_n1391_));
  NAND2_X1  g1026(.A1(new_n942_), .A2(new_n686_), .ZN(new_n1392_));
  NAND2_X1  g1027(.A1(new_n938_), .A2(new_n685_), .ZN(new_n1393_));
  OAI211_X1 g1028(.A(new_n1392_), .B(new_n1393_), .C1(new_n1374_), .C2(KEYINPUT53), .ZN(new_n1394_));
  XNOR2_X1  g1029(.A(new_n1394_), .B(new_n1375_), .ZN(new_n1395_));
  XNOR2_X1  g1030(.A(new_n1395_), .B(new_n677_), .ZN(new_n1396_));
  NOR2_X1   g1031(.A1(new_n1396_), .A2(new_n1390_), .ZN(new_n1397_));
  INV_X1    g1032(.A(new_n1397_), .ZN(new_n1398_));
  NAND2_X1  g1033(.A1(new_n1391_), .A2(new_n1398_), .ZN(new_n1399_));
  INV_X1    g1034(.A(new_n1399_), .ZN(new_n1400_));
  NAND2_X1  g1035(.A1(new_n1367_), .A2(new_n1400_), .ZN(new_n1401_));
  NAND3_X1  g1036(.A1(new_n1399_), .A2(new_n1341_), .A3(new_n1366_), .ZN(new_n1402_));
  NAND3_X1  g1037(.A1(new_n1401_), .A2(G4091), .A3(new_n1402_), .ZN(new_n1403_));
  INV_X1    g1038(.A(new_n1403_), .ZN(new_n1404_));
  NAND2_X1  g1039(.A1(new_n441_), .A2(new_n458_), .ZN(new_n1405_));
  NAND2_X1  g1040(.A1(new_n529_), .A2(G324), .ZN(new_n1406_));
  AOI21_X1  g1041(.A(G503), .B1(new_n1405_), .B2(new_n1406_), .ZN(new_n1407_));
  NAND2_X1  g1042(.A1(G248), .A2(G324), .ZN(new_n1408_));
  OAI21_X1  g1043(.A(new_n1408_), .B1(new_n429_), .B2(G324), .ZN(new_n1409_));
  AOI21_X1  g1044(.A(new_n1407_), .B1(G503), .B2(new_n1409_), .ZN(new_n1410_));
  NAND2_X1  g1045(.A1(G248), .A2(G514), .ZN(new_n1411_));
  OAI21_X1  g1046(.A(new_n1411_), .B1(G242), .B2(G514), .ZN(new_n1412_));
  XNOR2_X1  g1047(.A(new_n1410_), .B(new_n1412_), .ZN(new_n1413_));
  NAND2_X1  g1048(.A1(new_n441_), .A2(new_n637_), .ZN(new_n1414_));
  NAND2_X1  g1049(.A1(new_n529_), .A2(G341), .ZN(new_n1415_));
  AOI21_X1  g1050(.A(G523), .B1(new_n1414_), .B2(new_n1415_), .ZN(new_n1416_));
  OAI22_X1  g1051(.A1(new_n451_), .A2(new_n429_), .B1(new_n430_), .B2(new_n637_), .ZN(new_n1417_));
  AOI21_X1  g1052(.A(new_n1416_), .B1(new_n1417_), .B2(G523), .ZN(new_n1418_));
  XNOR2_X1  g1053(.A(new_n1413_), .B(new_n1418_), .ZN(new_n1419_));
  XNOR2_X1  g1054(.A(new_n432_), .B(new_n439_), .ZN(new_n1420_));
  XOR2_X1   g1055(.A(new_n445_), .B(new_n442_), .Z(new_n1421_));
  XNOR2_X1  g1056(.A(new_n1420_), .B(new_n1421_), .ZN(new_n1422_));
  XNOR2_X1  g1057(.A(new_n1419_), .B(new_n1422_), .ZN(new_n1423_));
  NOR2_X1   g1058(.A1(new_n468_), .A2(G242), .ZN(new_n1424_));
  NOR2_X1   g1059(.A1(G254), .A2(G351), .ZN(new_n1425_));
  OAI21_X1  g1060(.A(new_n624_), .B1(new_n1424_), .B2(new_n1425_), .ZN(new_n1426_));
  MUX2_X1   g1061(.A(new_n429_), .B(new_n430_), .S(G351), .Z(new_n1427_));
  OAI21_X1  g1062(.A(new_n1426_), .B1(new_n1427_), .B2(new_n624_), .ZN(new_n1428_));
  XNOR2_X1  g1063(.A(new_n1428_), .B(new_n752_), .ZN(new_n1429_));
  AND2_X1   g1064(.A1(new_n1423_), .A2(new_n1429_), .ZN(new_n1430_));
  OAI21_X1  g1065(.A(new_n753_), .B1(new_n1423_), .B2(new_n1429_), .ZN(new_n1431_));
  OAI21_X1  g1066(.A(new_n756_), .B1(new_n1430_), .B2(new_n1431_), .ZN(new_n1432_));
  OAI21_X1  g1067(.A(new_n1262_), .B1(new_n1404_), .B2(new_n1432_), .ZN(G843));
  NAND2_X1  g1068(.A1(new_n724_), .A2(new_n598_), .ZN(new_n1434_));
  NAND3_X1  g1069(.A1(new_n723_), .A2(new_n607_), .A3(new_n597_), .ZN(new_n1435_));
  NAND3_X1  g1070(.A1(new_n1434_), .A2(new_n619_), .A3(new_n1435_), .ZN(new_n1436_));
  OR2_X1    g1071(.A1(new_n1436_), .A2(KEYINPUT56), .ZN(new_n1437_));
  NAND2_X1  g1072(.A1(new_n1436_), .A2(KEYINPUT56), .ZN(new_n1438_));
  NAND2_X1  g1073(.A1(new_n1437_), .A2(new_n1438_), .ZN(new_n1439_));
  AOI21_X1  g1074(.A(new_n594_), .B1(new_n1434_), .B2(new_n1435_), .ZN(new_n1440_));
  AOI211_X1 g1075(.A(new_n509_), .B(new_n593_), .C1(new_n723_), .C2(new_n607_), .ZN(new_n1441_));
  OAI21_X1  g1076(.A(new_n616_), .B1(new_n1440_), .B2(new_n1441_), .ZN(new_n1442_));
  NOR2_X1   g1077(.A1(new_n1440_), .A2(new_n1441_), .ZN(new_n1443_));
  NAND2_X1  g1078(.A1(new_n1443_), .A2(new_n618_), .ZN(new_n1444_));
  NAND3_X1  g1079(.A1(new_n1439_), .A2(new_n1442_), .A3(new_n1444_), .ZN(new_n1445_));
  XNOR2_X1  g1080(.A(new_n604_), .B(new_n609_), .ZN(new_n1446_));
  OR2_X1    g1081(.A1(new_n1445_), .A2(new_n1446_), .ZN(new_n1447_));
  NAND2_X1  g1082(.A1(new_n1445_), .A2(new_n1446_), .ZN(new_n1448_));
  NAND2_X1  g1083(.A1(new_n734_), .A2(new_n590_), .ZN(new_n1449_));
  INV_X1    g1084(.A(G1497), .ZN(new_n1450_));
  NOR2_X1   g1085(.A1(new_n1449_), .A2(new_n1450_), .ZN(new_n1451_));
  NAND3_X1  g1086(.A1(new_n1447_), .A2(new_n1448_), .A3(new_n1451_), .ZN(new_n1452_));
  NAND2_X1  g1087(.A1(new_n1452_), .A2(KEYINPUT57), .ZN(new_n1453_));
  INV_X1    g1088(.A(KEYINPUT57), .ZN(new_n1454_));
  NAND4_X1  g1089(.A1(new_n1447_), .A2(new_n1454_), .A3(new_n1448_), .A4(new_n1451_), .ZN(new_n1455_));
  NAND2_X1  g1090(.A1(new_n1453_), .A2(new_n1455_), .ZN(new_n1456_));
  NOR2_X1   g1091(.A1(new_n596_), .A2(new_n617_), .ZN(new_n1457_));
  AOI21_X1  g1092(.A(new_n1457_), .B1(new_n596_), .B2(new_n616_), .ZN(new_n1458_));
  AND3_X1   g1093(.A1(new_n902_), .A2(new_n607_), .A3(new_n1458_), .ZN(new_n1459_));
  AOI21_X1  g1094(.A(new_n1458_), .B1(new_n902_), .B2(new_n607_), .ZN(new_n1460_));
  OR3_X1    g1095(.A1(new_n1459_), .A2(new_n1460_), .A3(new_n604_), .ZN(new_n1461_));
  OAI21_X1  g1096(.A(new_n604_), .B1(new_n1459_), .B2(new_n1460_), .ZN(new_n1462_));
  NAND2_X1  g1097(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1463_));
  XNOR2_X1  g1098(.A(new_n597_), .B(new_n619_), .ZN(new_n1464_));
  XNOR2_X1  g1099(.A(new_n1464_), .B(new_n609_), .ZN(new_n1465_));
  XNOR2_X1  g1100(.A(new_n1463_), .B(new_n1465_), .ZN(new_n1466_));
  AOI21_X1  g1101(.A(G1497), .B1(new_n1466_), .B2(new_n897_), .ZN(new_n1467_));
  AND2_X1   g1102(.A1(new_n1447_), .A2(new_n1448_), .ZN(new_n1468_));
  OAI21_X1  g1103(.A(new_n1467_), .B1(new_n1468_), .B2(new_n897_), .ZN(new_n1469_));
  AOI211_X1 g1104(.A(new_n1450_), .B(new_n1466_), .C1(new_n590_), .C2(new_n734_), .ZN(new_n1470_));
  INV_X1    g1105(.A(new_n1470_), .ZN(new_n1471_));
  NAND3_X1  g1106(.A1(new_n1456_), .A2(new_n1469_), .A3(new_n1471_), .ZN(new_n1472_));
  AOI21_X1  g1107(.A(new_n726_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n1473_));
  OAI21_X1  g1108(.A(new_n563_), .B1(new_n566_), .B2(new_n1473_), .ZN(new_n1474_));
  INV_X1    g1109(.A(KEYINPUT58), .ZN(new_n1475_));
  NAND2_X1  g1110(.A1(new_n1474_), .A2(new_n1475_), .ZN(new_n1476_));
  OAI211_X1 g1111(.A(KEYINPUT58), .B(new_n563_), .C1(new_n566_), .C2(new_n1473_), .ZN(new_n1477_));
  OAI211_X1 g1112(.A(new_n1476_), .B(new_n1477_), .C1(new_n564_), .C2(new_n730_), .ZN(new_n1478_));
  INV_X1    g1113(.A(new_n1478_), .ZN(new_n1479_));
  NOR2_X1   g1114(.A1(new_n863_), .A2(new_n726_), .ZN(new_n1480_));
  NAND2_X1  g1115(.A1(new_n1480_), .A2(new_n588_), .ZN(new_n1481_));
  INV_X1    g1116(.A(new_n1481_), .ZN(new_n1482_));
  OAI21_X1  g1117(.A(new_n730_), .B1(new_n1473_), .B2(new_n554_), .ZN(new_n1483_));
  NAND2_X1  g1118(.A1(new_n1483_), .A2(new_n770_), .ZN(new_n1484_));
  OAI211_X1 g1119(.A(new_n730_), .B(new_n587_), .C1(new_n1473_), .C2(new_n554_), .ZN(new_n1485_));
  NAND2_X1  g1120(.A1(new_n1484_), .A2(new_n1485_), .ZN(new_n1486_));
  NOR2_X1   g1121(.A1(new_n1482_), .A2(new_n1486_), .ZN(new_n1487_));
  AOI21_X1  g1122(.A(new_n1481_), .B1(new_n1484_), .B2(new_n1485_), .ZN(new_n1488_));
  OAI21_X1  g1123(.A(new_n1479_), .B1(new_n1487_), .B2(new_n1488_), .ZN(new_n1489_));
  AND2_X1   g1124(.A1(new_n1484_), .A2(new_n1485_), .ZN(new_n1490_));
  NAND3_X1  g1125(.A1(new_n1490_), .A2(KEYINPUT59), .A3(new_n1481_), .ZN(new_n1491_));
  INV_X1    g1126(.A(KEYINPUT59), .ZN(new_n1492_));
  OAI21_X1  g1127(.A(new_n1482_), .B1(new_n1486_), .B2(new_n1492_), .ZN(new_n1493_));
  NAND3_X1  g1128(.A1(new_n1491_), .A2(new_n1478_), .A3(new_n1493_), .ZN(new_n1494_));
  NAND2_X1  g1129(.A1(new_n1489_), .A2(new_n1494_), .ZN(new_n1495_));
  NAND2_X1  g1130(.A1(new_n1495_), .A2(new_n771_), .ZN(new_n1496_));
  INV_X1    g1131(.A(new_n771_), .ZN(new_n1497_));
  NAND3_X1  g1132(.A1(new_n1489_), .A2(new_n1494_), .A3(new_n1497_), .ZN(new_n1498_));
  NAND3_X1  g1133(.A1(new_n1496_), .A2(new_n840_), .A3(new_n1498_), .ZN(new_n1499_));
  NAND2_X1  g1134(.A1(new_n1490_), .A2(new_n1481_), .ZN(new_n1500_));
  NAND2_X1  g1135(.A1(new_n1482_), .A2(new_n1486_), .ZN(new_n1501_));
  NAND3_X1  g1136(.A1(new_n1500_), .A2(new_n1478_), .A3(new_n1501_), .ZN(new_n1502_));
  NAND2_X1  g1137(.A1(new_n1502_), .A2(new_n1497_), .ZN(new_n1503_));
  AOI21_X1  g1138(.A(new_n1478_), .B1(new_n1491_), .B2(new_n1493_), .ZN(new_n1504_));
  NOR2_X1   g1139(.A1(new_n1503_), .A2(new_n1504_), .ZN(new_n1505_));
  AOI21_X1  g1140(.A(new_n1497_), .B1(new_n1489_), .B2(new_n1494_), .ZN(new_n1506_));
  OAI21_X1  g1141(.A(new_n586_), .B1(new_n1505_), .B2(new_n1506_), .ZN(new_n1507_));
  AND3_X1   g1142(.A1(new_n1499_), .A2(new_n1507_), .A3(new_n574_), .ZN(new_n1508_));
  AOI21_X1  g1143(.A(new_n574_), .B1(new_n1499_), .B2(new_n1507_), .ZN(new_n1509_));
  OAI21_X1  g1144(.A(new_n556_), .B1(new_n1508_), .B2(new_n1509_), .ZN(new_n1510_));
  NAND2_X1  g1145(.A1(new_n1499_), .A2(new_n1507_), .ZN(new_n1511_));
  NAND2_X1  g1146(.A1(new_n1511_), .A2(new_n575_), .ZN(new_n1512_));
  AND3_X1   g1147(.A1(new_n1489_), .A2(new_n1494_), .A3(new_n1497_), .ZN(new_n1513_));
  OAI21_X1  g1148(.A(new_n586_), .B1(new_n1513_), .B2(new_n1506_), .ZN(new_n1514_));
  AND2_X1   g1149(.A1(new_n1491_), .A2(new_n1493_), .ZN(new_n1515_));
  OAI211_X1 g1150(.A(new_n1497_), .B(new_n1502_), .C1(new_n1515_), .C2(new_n1478_), .ZN(new_n1516_));
  NAND3_X1  g1151(.A1(new_n1496_), .A2(new_n1516_), .A3(new_n840_), .ZN(new_n1517_));
  NAND3_X1  g1152(.A1(new_n1514_), .A2(new_n1517_), .A3(new_n574_), .ZN(new_n1518_));
  NAND3_X1  g1153(.A1(new_n1512_), .A2(new_n725_), .A3(new_n1518_), .ZN(new_n1519_));
  AND3_X1   g1154(.A1(new_n1510_), .A2(new_n1519_), .A3(new_n564_), .ZN(new_n1520_));
  AND3_X1   g1155(.A1(new_n1514_), .A2(new_n1517_), .A3(new_n574_), .ZN(new_n1521_));
  OAI21_X1  g1156(.A(new_n556_), .B1(new_n1521_), .B2(new_n1509_), .ZN(new_n1522_));
  NAND3_X1  g1157(.A1(new_n1499_), .A2(new_n1507_), .A3(new_n574_), .ZN(new_n1523_));
  NAND3_X1  g1158(.A1(new_n1512_), .A2(new_n725_), .A3(new_n1523_), .ZN(new_n1524_));
  AOI21_X1  g1159(.A(new_n564_), .B1(new_n1522_), .B2(new_n1524_), .ZN(new_n1525_));
  OAI21_X1  g1160(.A(G1497), .B1(new_n1520_), .B2(new_n1525_), .ZN(new_n1526_));
  OAI21_X1  g1161(.A(new_n579_), .B1(new_n728_), .B2(new_n555_), .ZN(new_n1527_));
  AOI21_X1  g1162(.A(new_n554_), .B1(new_n1480_), .B2(new_n730_), .ZN(new_n1528_));
  OAI21_X1  g1163(.A(new_n1527_), .B1(new_n1528_), .B2(new_n579_), .ZN(new_n1529_));
  XNOR2_X1  g1164(.A(new_n1529_), .B(new_n1497_), .ZN(new_n1530_));
  INV_X1    g1165(.A(new_n1480_), .ZN(new_n1531_));
  AOI21_X1  g1166(.A(new_n1531_), .B1(new_n732_), .B2(new_n563_), .ZN(new_n1532_));
  INV_X1    g1167(.A(new_n1532_), .ZN(new_n1533_));
  NAND3_X1  g1168(.A1(new_n732_), .A2(new_n563_), .A3(new_n1531_), .ZN(new_n1534_));
  AOI21_X1  g1169(.A(new_n586_), .B1(new_n1533_), .B2(new_n1534_), .ZN(new_n1535_));
  INV_X1    g1170(.A(new_n1535_), .ZN(new_n1536_));
  NAND3_X1  g1171(.A1(new_n1533_), .A2(new_n586_), .A3(new_n1534_), .ZN(new_n1537_));
  NAND3_X1  g1172(.A1(new_n1530_), .A2(new_n1536_), .A3(new_n1537_), .ZN(new_n1538_));
  XNOR2_X1  g1173(.A(new_n1529_), .B(new_n771_), .ZN(new_n1539_));
  INV_X1    g1174(.A(new_n1537_), .ZN(new_n1540_));
  OAI21_X1  g1175(.A(new_n1539_), .B1(new_n1540_), .B2(new_n1535_), .ZN(new_n1541_));
  NAND3_X1  g1176(.A1(new_n1538_), .A2(new_n1541_), .A3(new_n574_), .ZN(new_n1542_));
  AND2_X1   g1177(.A1(new_n725_), .A2(KEYINPUT60), .ZN(new_n1543_));
  NAND2_X1  g1178(.A1(new_n1542_), .A2(new_n1543_), .ZN(new_n1544_));
  AOI21_X1  g1179(.A(new_n574_), .B1(new_n1538_), .B2(new_n1541_), .ZN(new_n1545_));
  NAND2_X1  g1180(.A1(new_n1544_), .A2(new_n1545_), .ZN(new_n1546_));
  NAND2_X1  g1181(.A1(new_n1538_), .A2(new_n1541_), .ZN(new_n1547_));
  NAND2_X1  g1182(.A1(new_n1547_), .A2(new_n575_), .ZN(new_n1548_));
  NAND3_X1  g1183(.A1(new_n1548_), .A2(new_n1542_), .A3(new_n1543_), .ZN(new_n1549_));
  OR2_X1    g1184(.A1(new_n1542_), .A2(new_n725_), .ZN(new_n1550_));
  NAND4_X1  g1185(.A1(new_n1546_), .A2(new_n1549_), .A3(new_n564_), .A4(new_n1550_), .ZN(new_n1551_));
  NAND2_X1  g1186(.A1(new_n1551_), .A2(new_n1450_), .ZN(new_n1552_));
  NOR2_X1   g1187(.A1(new_n1542_), .A2(new_n725_), .ZN(new_n1553_));
  AOI21_X1  g1188(.A(new_n1553_), .B1(new_n1545_), .B2(new_n1544_), .ZN(new_n1554_));
  AOI21_X1  g1189(.A(new_n564_), .B1(new_n1554_), .B2(new_n1549_), .ZN(new_n1555_));
  OR2_X1    g1190(.A1(new_n1552_), .A2(new_n1555_), .ZN(new_n1556_));
  AOI21_X1  g1191(.A(new_n1472_), .B1(new_n1526_), .B2(new_n1556_), .ZN(new_n1557_));
  NOR3_X1   g1192(.A1(new_n1508_), .A2(new_n1509_), .A3(new_n556_), .ZN(new_n1558_));
  AOI21_X1  g1193(.A(new_n725_), .B1(new_n1512_), .B2(new_n1518_), .ZN(new_n1559_));
  OAI21_X1  g1194(.A(new_n565_), .B1(new_n1558_), .B2(new_n1559_), .ZN(new_n1560_));
  NAND3_X1  g1195(.A1(new_n1522_), .A2(new_n1524_), .A3(new_n564_), .ZN(new_n1561_));
  AOI21_X1  g1196(.A(new_n1450_), .B1(new_n1560_), .B2(new_n1561_), .ZN(new_n1562_));
  OAI21_X1  g1197(.A(new_n1472_), .B1(new_n1552_), .B2(new_n1555_), .ZN(new_n1563_));
  NOR2_X1   g1198(.A1(new_n1562_), .A2(new_n1563_), .ZN(new_n1564_));
  OAI21_X1  g1199(.A(new_n762_), .B1(new_n1557_), .B2(new_n1564_), .ZN(new_n1565_));
  OAI21_X1  g1200(.A(G4092), .B1(G118), .B2(G4091), .ZN(new_n1566_));
  NOR2_X1   g1201(.A1(new_n479_), .A2(G242), .ZN(new_n1567_));
  NOR2_X1   g1202(.A1(G218), .A2(G254), .ZN(new_n1568_));
  OAI21_X1  g1203(.A(new_n614_), .B1(new_n1567_), .B2(new_n1568_), .ZN(new_n1569_));
  MUX2_X1   g1204(.A(new_n429_), .B(new_n430_), .S(G218), .Z(new_n1570_));
  OAI21_X1  g1205(.A(new_n1569_), .B1(new_n1570_), .B2(new_n614_), .ZN(new_n1571_));
  NOR2_X1   g1206(.A1(new_n510_), .A2(G242), .ZN(new_n1572_));
  NOR2_X1   g1207(.A1(G226), .A2(G254), .ZN(new_n1573_));
  OAI21_X1  g1208(.A(new_n509_), .B1(new_n1572_), .B2(new_n1573_), .ZN(new_n1574_));
  MUX2_X1   g1209(.A(new_n429_), .B(new_n430_), .S(G226), .Z(new_n1575_));
  OAI21_X1  g1210(.A(new_n1574_), .B1(new_n1575_), .B2(new_n509_), .ZN(new_n1576_));
  XNOR2_X1  g1211(.A(new_n1571_), .B(new_n1576_), .ZN(new_n1577_));
  XNOR2_X1  g1212(.A(new_n1577_), .B(new_n536_), .ZN(new_n1578_));
  NAND2_X1  g1213(.A1(new_n496_), .A2(new_n441_), .ZN(new_n1579_));
  NAND2_X1  g1214(.A1(new_n529_), .A2(G210), .ZN(new_n1580_));
  AOI21_X1  g1215(.A(G457), .B1(new_n1579_), .B2(new_n1580_), .ZN(new_n1581_));
  NAND2_X1  g1216(.A1(G210), .A2(G248), .ZN(new_n1582_));
  OAI21_X1  g1217(.A(new_n1582_), .B1(new_n429_), .B2(G210), .ZN(new_n1583_));
  AOI21_X1  g1218(.A(new_n1581_), .B1(G457), .B2(new_n1583_), .ZN(new_n1584_));
  XNOR2_X1  g1219(.A(new_n1578_), .B(new_n1584_), .ZN(new_n1585_));
  OAI21_X1  g1220(.A(new_n561_), .B1(new_n529_), .B2(new_n490_), .ZN(new_n1586_));
  AOI22_X1  g1221(.A1(new_n1586_), .A2(KEYINPUT61), .B1(G254), .B2(new_n490_), .ZN(new_n1587_));
  OAI21_X1  g1222(.A(new_n1587_), .B1(KEYINPUT61), .B2(new_n1586_), .ZN(new_n1588_));
  NOR2_X1   g1223(.A1(new_n430_), .A2(new_n490_), .ZN(new_n1589_));
  NOR2_X1   g1224(.A1(new_n429_), .A2(G257), .ZN(new_n1590_));
  OAI21_X1  g1225(.A(G389), .B1(new_n1589_), .B2(new_n1590_), .ZN(new_n1591_));
  NAND2_X1  g1226(.A1(new_n1588_), .A2(new_n1591_), .ZN(new_n1592_));
  NOR2_X1   g1227(.A1(new_n505_), .A2(G242), .ZN(new_n1593_));
  NOR2_X1   g1228(.A1(G234), .A2(G254), .ZN(new_n1594_));
  OAI21_X1  g1229(.A(new_n570_), .B1(new_n1593_), .B2(new_n1594_), .ZN(new_n1595_));
  MUX2_X1   g1230(.A(new_n429_), .B(new_n430_), .S(G234), .Z(new_n1596_));
  OAI21_X1  g1231(.A(new_n1595_), .B1(new_n1596_), .B2(new_n570_), .ZN(new_n1597_));
  XNOR2_X1  g1232(.A(new_n1592_), .B(new_n1597_), .ZN(new_n1598_));
  XNOR2_X1  g1233(.A(new_n1585_), .B(new_n1598_), .ZN(new_n1599_));
  NOR2_X1   g1234(.A1(new_n519_), .A2(G242), .ZN(new_n1600_));
  NOR2_X1   g1235(.A1(G254), .A2(G273), .ZN(new_n1601_));
  OAI21_X1  g1236(.A(new_n518_), .B1(new_n1600_), .B2(new_n1601_), .ZN(new_n1602_));
  MUX2_X1   g1237(.A(new_n429_), .B(new_n430_), .S(G273), .Z(new_n1603_));
  OAI21_X1  g1238(.A(new_n1602_), .B1(new_n1603_), .B2(new_n518_), .ZN(new_n1604_));
  NOR2_X1   g1239(.A1(new_n484_), .A2(G242), .ZN(new_n1605_));
  NOR2_X1   g1240(.A1(G254), .A2(G265), .ZN(new_n1606_));
  OAI21_X1  g1241(.A(new_n552_), .B1(new_n1605_), .B2(new_n1606_), .ZN(new_n1607_));
  MUX2_X1   g1242(.A(new_n429_), .B(new_n430_), .S(G265), .Z(new_n1608_));
  OAI21_X1  g1243(.A(new_n1607_), .B1(new_n1608_), .B2(new_n552_), .ZN(new_n1609_));
  XNOR2_X1  g1244(.A(new_n1604_), .B(new_n1609_), .ZN(new_n1610_));
  NAND2_X1  g1245(.A1(new_n441_), .A2(new_n538_), .ZN(new_n1611_));
  NAND2_X1  g1246(.A1(new_n529_), .A2(G281), .ZN(new_n1612_));
  AOI21_X1  g1247(.A(G374), .B1(new_n1611_), .B2(new_n1612_), .ZN(new_n1613_));
  NAND2_X1  g1248(.A1(G248), .A2(G281), .ZN(new_n1614_));
  OAI21_X1  g1249(.A(new_n1614_), .B1(new_n429_), .B2(G281), .ZN(new_n1615_));
  AOI21_X1  g1250(.A(new_n1613_), .B1(G374), .B2(new_n1615_), .ZN(new_n1616_));
  XNOR2_X1  g1251(.A(new_n1610_), .B(new_n1616_), .ZN(new_n1617_));
  XNOR2_X1  g1252(.A(new_n1599_), .B(new_n1617_), .ZN(new_n1618_));
  NAND3_X1  g1253(.A1(new_n1618_), .A2(new_n753_), .A3(new_n756_), .ZN(new_n1619_));
  XNOR2_X1  g1254(.A(new_n1619_), .B(KEYINPUT62), .ZN(new_n1620_));
  NAND3_X1  g1255(.A1(new_n1565_), .A2(new_n1566_), .A3(new_n1620_), .ZN(G882));
  NAND2_X1  g1256(.A1(G64), .A2(G4088), .ZN(new_n1622_));
  INV_X1    g1257(.A(G14), .ZN(new_n1623_));
  OAI21_X1  g1258(.A(new_n1622_), .B1(new_n1623_), .B2(G4088), .ZN(new_n1624_));
  NAND2_X1  g1259(.A1(new_n1624_), .A2(G4087), .ZN(new_n1625_));
  NAND2_X1  g1260(.A1(new_n1618_), .A2(new_n753_), .ZN(new_n1626_));
  NAND2_X1  g1261(.A1(new_n1626_), .A2(new_n756_), .ZN(new_n1627_));
  INV_X1    g1262(.A(new_n1627_), .ZN(new_n1628_));
  NAND2_X1  g1263(.A1(new_n1565_), .A2(new_n1628_), .ZN(new_n1629_));
  NAND2_X1  g1264(.A1(G97), .A2(G4092), .ZN(new_n1630_));
  AOI21_X1  g1265(.A(new_n787_), .B1(new_n1629_), .B2(new_n1630_), .ZN(new_n1631_));
  NAND2_X1  g1266(.A1(G94), .A2(G4092), .ZN(new_n1632_));
  NOR2_X1   g1267(.A1(new_n1430_), .A2(new_n1431_), .ZN(new_n1633_));
  XNOR2_X1  g1268(.A(new_n1633_), .B(KEYINPUT63), .ZN(new_n1634_));
  INV_X1    g1269(.A(new_n1634_), .ZN(new_n1635_));
  AOI21_X1  g1270(.A(new_n753_), .B1(new_n1367_), .B2(new_n1400_), .ZN(new_n1636_));
  AOI21_X1  g1271(.A(new_n1635_), .B1(new_n1636_), .B2(new_n1402_), .ZN(new_n1637_));
  OAI21_X1  g1272(.A(new_n1632_), .B1(new_n1637_), .B2(G4092), .ZN(new_n1638_));
  AOI21_X1  g1273(.A(new_n1631_), .B1(new_n787_), .B2(new_n1638_), .ZN(new_n1639_));
  OAI21_X1  g1274(.A(new_n1625_), .B1(new_n1639_), .B2(G4087), .ZN(G767));
  NAND2_X1  g1275(.A1(G64), .A2(G4089), .ZN(new_n1641_));
  OAI21_X1  g1276(.A(new_n1641_), .B1(new_n1623_), .B2(G4089), .ZN(new_n1642_));
  NAND2_X1  g1277(.A1(new_n1642_), .A2(G4090), .ZN(new_n1643_));
  AOI21_X1  g1278(.A(new_n830_), .B1(new_n1629_), .B2(new_n1630_), .ZN(new_n1644_));
  AOI21_X1  g1279(.A(new_n1644_), .B1(new_n830_), .B2(new_n1638_), .ZN(new_n1645_));
  OAI21_X1  g1280(.A(new_n1643_), .B1(new_n1645_), .B2(G4090), .ZN(G807));
  AOI21_X1  g1281(.A(G4092), .B1(new_n1403_), .B2(new_n1634_), .ZN(new_n1647_));
  INV_X1    g1282(.A(new_n1632_), .ZN(new_n1648_));
  OAI21_X1  g1283(.A(new_n954_), .B1(new_n1647_), .B2(new_n1648_), .ZN(new_n1649_));
  INV_X1    g1284(.A(new_n1472_), .ZN(new_n1650_));
  NAND3_X1  g1285(.A1(new_n1510_), .A2(new_n1519_), .A3(new_n564_), .ZN(new_n1651_));
  AOI21_X1  g1286(.A(new_n1450_), .B1(new_n1560_), .B2(new_n1651_), .ZN(new_n1652_));
  NOR2_X1   g1287(.A1(new_n1552_), .A2(new_n1555_), .ZN(new_n1653_));
  OAI21_X1  g1288(.A(new_n1650_), .B1(new_n1652_), .B2(new_n1653_), .ZN(new_n1654_));
  INV_X1    g1289(.A(new_n1561_), .ZN(new_n1655_));
  OAI21_X1  g1290(.A(G1497), .B1(new_n1655_), .B2(new_n1525_), .ZN(new_n1656_));
  NAND3_X1  g1291(.A1(new_n1656_), .A2(new_n1556_), .A3(new_n1472_), .ZN(new_n1657_));
  AOI21_X1  g1292(.A(new_n763_), .B1(new_n1654_), .B2(new_n1657_), .ZN(new_n1658_));
  OAI21_X1  g1293(.A(new_n1630_), .B1(new_n1658_), .B2(new_n1627_), .ZN(new_n1659_));
  NAND2_X1  g1294(.A1(new_n1659_), .A2(G1689), .ZN(new_n1660_));
  AOI21_X1  g1295(.A(G1690), .B1(new_n1649_), .B2(new_n1660_), .ZN(new_n1661_));
  NAND2_X1  g1296(.A1(new_n954_), .A2(G176), .ZN(new_n1662_));
  NAND2_X1  g1297(.A1(G179), .A2(G1689), .ZN(new_n1663_));
  AOI21_X1  g1298(.A(new_n953_), .B1(new_n1662_), .B2(new_n1663_), .ZN(new_n1664_));
  OAI21_X1  g1299(.A(G137), .B1(new_n1661_), .B2(new_n1664_), .ZN(G658));
  OAI21_X1  g1300(.A(new_n1069_), .B1(new_n1647_), .B2(new_n1648_), .ZN(new_n1666_));
  NAND2_X1  g1301(.A1(new_n1659_), .A2(G1691), .ZN(new_n1667_));
  AOI21_X1  g1302(.A(G1694), .B1(new_n1666_), .B2(new_n1667_), .ZN(new_n1668_));
  NAND2_X1  g1303(.A1(new_n1069_), .A2(G176), .ZN(new_n1669_));
  NAND2_X1  g1304(.A1(G179), .A2(G1691), .ZN(new_n1670_));
  AOI21_X1  g1305(.A(new_n966_), .B1(new_n1669_), .B2(new_n1670_), .ZN(new_n1671_));
  OAI21_X1  g1306(.A(G137), .B1(new_n1668_), .B2(new_n1671_), .ZN(G690));
endmodule


