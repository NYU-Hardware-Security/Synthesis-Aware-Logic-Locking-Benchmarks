//Secret key is'0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_c1355" written by ABC on Tue Nov  1 15:33:44 2022

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n460_, new_n461_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n492_, new_n493_, new_n494_, new_n496_, new_n497_, new_n498_,
    new_n500_, new_n501_, new_n502_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n520_,
    new_n521_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n601_, new_n603_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_;
  INV_X1    g000(.A(G127gat), .ZN(new_n138_));
  NOR2_X1   g001(.A1(new_n138_), .A2(G134gat), .ZN(new_n139_));
  INV_X1    g002(.A(G134gat), .ZN(new_n140_));
  NOR2_X1   g003(.A1(new_n140_), .A2(G127gat), .ZN(new_n141_));
  OAI21_X1  g004(.A(KEYINPUT1), .B1(new_n139_), .B2(new_n141_), .ZN(new_n142_));
  NAND2_X1  g005(.A1(new_n140_), .A2(G127gat), .ZN(new_n143_));
  NAND2_X1  g006(.A1(new_n138_), .A2(G134gat), .ZN(new_n144_));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n145_));
  NAND3_X1  g008(.A1(new_n143_), .A2(new_n144_), .A3(new_n145_), .ZN(new_n146_));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n147_));
  NAND3_X1  g010(.A1(new_n142_), .A2(new_n146_), .A3(new_n147_), .ZN(new_n148_));
  INV_X1    g011(.A(KEYINPUT4), .ZN(new_n149_));
  INV_X1    g012(.A(new_n147_), .ZN(new_n150_));
  NAND2_X1  g013(.A1(new_n143_), .A2(new_n144_), .ZN(new_n151_));
  NAND3_X1  g014(.A1(new_n150_), .A2(KEYINPUT1), .A3(new_n151_), .ZN(new_n152_));
  AND3_X1   g015(.A1(new_n148_), .A2(new_n149_), .A3(new_n152_), .ZN(new_n153_));
  AOI21_X1  g016(.A(new_n149_), .B1(new_n148_), .B2(new_n152_), .ZN(new_n154_));
  NOR2_X1   g017(.A1(new_n153_), .A2(new_n154_), .ZN(new_n155_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n156_));
  NAND2_X1  g019(.A1(new_n156_), .A2(KEYINPUT25), .ZN(new_n157_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n158_));
  NAND3_X1  g021(.A1(new_n158_), .A2(G183gat), .A3(G190gat), .ZN(new_n159_));
  OR2_X1    g022(.A1(G183gat), .A2(G190gat), .ZN(new_n160_));
  NAND3_X1  g023(.A1(new_n157_), .A2(new_n159_), .A3(new_n160_), .ZN(new_n161_));
  INV_X1    g024(.A(G169gat), .ZN(new_n162_));
  INV_X1    g025(.A(G176gat), .ZN(new_n163_));
  NAND3_X1  g026(.A1(new_n162_), .A2(new_n163_), .A3(KEYINPUT24), .ZN(new_n164_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n165_));
  OAI21_X1  g028(.A(new_n165_), .B1(G169gat), .B2(G176gat), .ZN(new_n166_));
  NAND2_X1  g029(.A1(new_n164_), .A2(new_n166_), .ZN(new_n167_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n168_));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n169_));
  NAND2_X1  g032(.A1(new_n168_), .A2(new_n169_), .ZN(new_n170_));
  NAND3_X1  g033(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n171_));
  NAND2_X1  g034(.A1(new_n170_), .A2(new_n171_), .ZN(new_n172_));
  NAND3_X1  g035(.A1(new_n161_), .A2(new_n167_), .A3(new_n172_), .ZN(new_n173_));
  INV_X1    g036(.A(G183gat), .ZN(new_n174_));
  AND2_X1   g037(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n175_));
  NOR2_X1   g038(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n176_));
  OAI21_X1  g039(.A(new_n174_), .B1(new_n175_), .B2(new_n176_), .ZN(new_n177_));
  XNOR2_X1  g040(.A(G169gat), .B(G176gat), .ZN(new_n178_));
  NAND3_X1  g041(.A1(new_n177_), .A2(new_n178_), .A3(new_n156_), .ZN(new_n179_));
  NAND2_X1  g042(.A1(new_n173_), .A2(new_n179_), .ZN(new_n180_));
  XOR2_X1   g043(.A(new_n155_), .B(new_n180_), .Z(new_n181_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n182_));
  XNOR2_X1  g045(.A(new_n181_), .B(new_n182_), .ZN(new_n183_));
  INV_X1    g046(.A(KEYINPUT31), .ZN(new_n184_));
  NAND2_X1  g047(.A1(new_n183_), .A2(new_n184_), .ZN(new_n185_));
  XNOR2_X1  g048(.A(G15gat), .B(G43gat), .ZN(new_n186_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n187_));
  XNOR2_X1  g050(.A(new_n186_), .B(new_n187_), .ZN(new_n188_));
  NAND2_X1  g051(.A1(new_n185_), .A2(new_n188_), .ZN(new_n189_));
  INV_X1    g052(.A(new_n188_), .ZN(new_n190_));
  NAND3_X1  g053(.A1(new_n183_), .A2(new_n184_), .A3(new_n190_), .ZN(new_n191_));
  NAND2_X1  g054(.A1(new_n189_), .A2(new_n191_), .ZN(new_n192_));
  INV_X1    g055(.A(G155gat), .ZN(new_n193_));
  INV_X1    g056(.A(G162gat), .ZN(new_n194_));
  NAND2_X1  g057(.A1(new_n193_), .A2(new_n194_), .ZN(new_n195_));
  INV_X1    g058(.A(G148gat), .ZN(new_n196_));
  NAND2_X1  g059(.A1(new_n196_), .A2(G141gat), .ZN(new_n197_));
  INV_X1    g060(.A(G141gat), .ZN(new_n198_));
  NAND2_X1  g061(.A1(new_n198_), .A2(G148gat), .ZN(new_n199_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n200_));
  NAND4_X1  g063(.A1(new_n195_), .A2(new_n197_), .A3(new_n199_), .A4(new_n200_), .ZN(new_n201_));
  NAND2_X1  g064(.A1(new_n201_), .A2(KEYINPUT3), .ZN(new_n202_));
  XNOR2_X1  g065(.A(G141gat), .B(G148gat), .ZN(new_n203_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n204_));
  NAND4_X1  g067(.A1(new_n203_), .A2(new_n204_), .A3(new_n200_), .A4(new_n195_), .ZN(new_n205_));
  OAI21_X1  g068(.A(KEYINPUT2), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  INV_X1    g069(.A(new_n206_), .ZN(new_n207_));
  NOR3_X1   g070(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n208_));
  OAI21_X1  g071(.A(new_n200_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g072(.A(new_n203_), .ZN(new_n210_));
  AOI22_X1  g073(.A1(new_n202_), .A2(new_n205_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g074(.A(G197gat), .B(G204gat), .Z(new_n212_));
  NOR2_X1   g075(.A1(G211gat), .A2(G218gat), .ZN(new_n213_));
  NAND2_X1  g076(.A1(G211gat), .A2(G218gat), .ZN(new_n214_));
  AOI21_X1  g077(.A(new_n213_), .B1(KEYINPUT21), .B2(new_n214_), .ZN(new_n215_));
  AND2_X1   g078(.A1(new_n213_), .A2(KEYINPUT21), .ZN(new_n216_));
  OAI21_X1  g079(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g080(.A(G211gat), .ZN(new_n218_));
  AND2_X1   g081(.A1(KEYINPUT22), .A2(G218gat), .ZN(new_n219_));
  NOR2_X1   g082(.A1(KEYINPUT22), .A2(G218gat), .ZN(new_n220_));
  OAI21_X1  g083(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n222_));
  NAND3_X1  g085(.A1(new_n221_), .A2(new_n214_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g086(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g087(.A(new_n211_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g088(.A(G228gat), .ZN(new_n226_));
  INV_X1    g089(.A(G233gat), .ZN(new_n227_));
  OAI21_X1  g090(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n229_));
  NAND2_X1  g092(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n231_));
  XNOR2_X1  g094(.A(new_n231_), .B(KEYINPUT29), .ZN(new_n232_));
  XOR2_X1   g095(.A(G22gat), .B(G50gat), .Z(new_n233_));
  XNOR2_X1  g096(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g097(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  OR3_X1    g098(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n236_));
  NAND2_X1  g099(.A1(new_n236_), .A2(new_n228_), .ZN(new_n237_));
  XNOR2_X1  g100(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g101(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g102(.A1(new_n192_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g103(.A(new_n211_), .ZN(new_n241_));
  OAI21_X1  g104(.A(new_n241_), .B1(new_n153_), .B2(new_n154_), .ZN(new_n242_));
  NAND2_X1  g105(.A1(new_n148_), .A2(new_n152_), .ZN(new_n243_));
  NAND2_X1  g106(.A1(new_n211_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  NAND3_X1  g108(.A1(new_n242_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  XOR2_X1   g109(.A(new_n245_), .B(KEYINPUT0), .Z(new_n247_));
  INV_X1    g110(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g111(.A(new_n244_), .ZN(new_n249_));
  NOR2_X1   g112(.A1(new_n211_), .A2(new_n243_), .ZN(new_n250_));
  OAI21_X1  g113(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n252_));
  XNOR2_X1  g115(.A(new_n252_), .B(G57gat), .ZN(new_n253_));
  INV_X1    g116(.A(G85gat), .ZN(new_n254_));
  XNOR2_X1  g117(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND3_X1  g118(.A1(new_n246_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g119(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g120(.A(new_n255_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n258_));
  NOR2_X1   g121(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g122(.A(new_n259_), .ZN(new_n260_));
  AND2_X1   g123(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  NAND4_X1  g124(.A1(new_n217_), .A2(new_n173_), .A3(new_n179_), .A4(new_n223_), .ZN(new_n262_));
  AOI21_X1  g125(.A(new_n261_), .B1(new_n262_), .B2(KEYINPUT27), .ZN(new_n263_));
  NAND2_X1  g126(.A1(new_n224_), .A2(new_n180_), .ZN(new_n264_));
  NAND2_X1  g127(.A1(new_n264_), .A2(new_n262_), .ZN(new_n265_));
  NAND2_X1  g128(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g129(.A(new_n264_), .B(new_n262_), .C1(KEYINPUT27), .C2(new_n261_), .ZN(new_n267_));
  NAND2_X1  g130(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n269_));
  INV_X1    g132(.A(G64gat), .ZN(new_n270_));
  OR2_X1    g133(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g134(.A1(new_n269_), .A2(new_n270_), .ZN(new_n272_));
  NAND2_X1  g135(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g136(.A(G92gat), .ZN(new_n274_));
  NAND2_X1  g137(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g138(.A1(new_n271_), .A2(G92gat), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g139(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g140(.A1(new_n277_), .A2(KEYINPUT20), .ZN(new_n278_));
  INV_X1    g141(.A(KEYINPUT20), .ZN(new_n279_));
  NAND3_X1  g142(.A1(new_n275_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n280_));
  NAND2_X1  g143(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NOR3_X1   g144(.A1(new_n268_), .A2(new_n281_), .A3(KEYINPUT28), .ZN(new_n282_));
  AOI22_X1  g145(.A1(new_n266_), .A2(new_n267_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n283_));
  NOR2_X1   g146(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g147(.A(KEYINPUT28), .B1(new_n268_), .B2(new_n281_), .ZN(new_n285_));
  NAND2_X1  g148(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR3_X1   g149(.A1(new_n240_), .A2(new_n260_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g150(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g151(.A(KEYINPUT35), .ZN(new_n289_));
  AOI21_X1  g152(.A(new_n245_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n290_));
  NOR3_X1   g153(.A1(new_n249_), .A2(new_n250_), .A3(new_n248_), .ZN(new_n291_));
  NOR2_X1   g154(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g155(.A(new_n256_), .B1(new_n292_), .B2(new_n255_), .ZN(new_n293_));
  AOI21_X1  g156(.A(new_n293_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n294_));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n295_));
  AND3_X1   g158(.A1(new_n266_), .A2(new_n295_), .A3(new_n267_), .ZN(new_n296_));
  AOI21_X1  g159(.A(new_n295_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n297_));
  OAI21_X1  g160(.A(new_n277_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g161(.A(KEYINPUT34), .ZN(new_n299_));
  NAND2_X1  g162(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g163(.A(KEYINPUT34), .B(new_n277_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n301_));
  AOI21_X1  g164(.A(new_n259_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g165(.A(new_n283_), .ZN(new_n303_));
  AOI21_X1  g166(.A(new_n294_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g167(.A(new_n289_), .B1(new_n304_), .B2(new_n238_), .ZN(new_n305_));
  NOR2_X1   g168(.A1(new_n286_), .A2(new_n260_), .ZN(new_n306_));
  NAND2_X1  g169(.A1(new_n306_), .A2(new_n238_), .ZN(new_n307_));
  AOI211_X1 g170(.A(new_n283_), .B(new_n259_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n308_));
  OAI211_X1 g171(.A(KEYINPUT35), .B(new_n239_), .C1(new_n308_), .C2(new_n294_), .ZN(new_n309_));
  NAND3_X1  g172(.A1(new_n305_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g173(.A(KEYINPUT32), .ZN(new_n311_));
  AND3_X1   g174(.A1(new_n189_), .A2(new_n311_), .A3(new_n191_), .ZN(new_n312_));
  AOI21_X1  g175(.A(new_n311_), .B1(new_n189_), .B2(new_n191_), .ZN(new_n313_));
  NOR2_X1   g176(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AND3_X1   g177(.A1(new_n310_), .A2(KEYINPUT36), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g178(.A(KEYINPUT36), .B1(new_n310_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g179(.A(new_n288_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g180(.A(G43gat), .B(G50gat), .ZN(new_n318_));
  INV_X1    g181(.A(G29gat), .ZN(new_n319_));
  NAND2_X1  g182(.A1(new_n319_), .A2(KEYINPUT15), .ZN(new_n320_));
  XNOR2_X1  g183(.A(new_n318_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g184(.A(G36gat), .ZN(new_n322_));
  OAI21_X1  g185(.A(new_n322_), .B1(new_n319_), .B2(KEYINPUT15), .ZN(new_n323_));
  XOR2_X1   g186(.A(new_n321_), .B(new_n323_), .Z(new_n324_));
  XNOR2_X1  g187(.A(G1gat), .B(G8gat), .ZN(new_n325_));
  INV_X1    g188(.A(G15gat), .ZN(new_n326_));
  INV_X1    g189(.A(G22gat), .ZN(new_n327_));
  NOR2_X1   g190(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g191(.A(new_n325_), .B1(KEYINPUT16), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g192(.A(G15gat), .B(G22gat), .ZN(new_n330_));
  XNOR2_X1  g193(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  OR2_X1    g194(.A1(new_n324_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g195(.A1(new_n324_), .A2(new_n331_), .ZN(new_n333_));
  AND2_X1   g196(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g197(.A1(G229gat), .A2(G233gat), .ZN(new_n335_));
  NAND2_X1  g198(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g199(.A1(new_n332_), .A2(KEYINPUT17), .A3(new_n333_), .ZN(new_n337_));
  OR2_X1    g200(.A1(new_n333_), .A2(KEYINPUT17), .ZN(new_n338_));
  XNOR2_X1  g201(.A(new_n335_), .B(KEYINPUT14), .ZN(new_n339_));
  NAND3_X1  g202(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g203(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g204(.A(G113gat), .B(G141gat), .ZN(new_n342_));
  XNOR2_X1  g205(.A(new_n342_), .B(G169gat), .ZN(new_n343_));
  XOR2_X1   g206(.A(new_n343_), .B(G197gat), .Z(new_n344_));
  INV_X1    g207(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g208(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g209(.A1(new_n336_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n347_));
  NAND2_X1  g210(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g211(.A(G99gat), .ZN(new_n349_));
  INV_X1    g212(.A(G106gat), .ZN(new_n350_));
  NAND2_X1  g213(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g214(.A1(G99gat), .A2(G106gat), .ZN(new_n352_));
  NOR2_X1   g215(.A1(new_n254_), .A2(new_n274_), .ZN(new_n353_));
  NOR2_X1   g216(.A1(G85gat), .A2(G92gat), .ZN(new_n354_));
  OAI211_X1 g217(.A(new_n351_), .B(new_n352_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g218(.A(new_n355_), .B(KEYINPUT9), .ZN(new_n356_));
  NAND2_X1  g219(.A1(new_n351_), .A2(KEYINPUT8), .ZN(new_n357_));
  INV_X1    g220(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g221(.A1(new_n351_), .A2(KEYINPUT8), .ZN(new_n359_));
  OAI21_X1  g222(.A(new_n352_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g223(.A(KEYINPUT7), .ZN(new_n361_));
  NAND2_X1  g224(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g225(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n363_));
  AOI21_X1  g226(.A(new_n353_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g227(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g228(.A1(new_n356_), .A2(new_n365_), .ZN(new_n366_));
  AND2_X1   g229(.A1(new_n366_), .A2(KEYINPUT11), .ZN(new_n367_));
  NOR2_X1   g230(.A1(new_n366_), .A2(KEYINPUT11), .ZN(new_n368_));
  OAI21_X1  g231(.A(new_n324_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g232(.A1(new_n369_), .A2(KEYINPUT37), .ZN(new_n370_));
  OR2_X1    g233(.A1(new_n324_), .A2(new_n366_), .ZN(new_n371_));
  XNOR2_X1  g234(.A(new_n366_), .B(KEYINPUT11), .ZN(new_n372_));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n373_));
  NAND3_X1  g236(.A1(new_n372_), .A2(new_n373_), .A3(new_n324_), .ZN(new_n374_));
  NAND3_X1  g237(.A1(new_n370_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g238(.A1(new_n375_), .A2(G232gat), .A3(G233gat), .ZN(new_n376_));
  INV_X1    g239(.A(G218gat), .ZN(new_n377_));
  NAND2_X1  g240(.A1(G232gat), .A2(G233gat), .ZN(new_n378_));
  NAND4_X1  g241(.A1(new_n370_), .A2(new_n374_), .A3(new_n378_), .A4(new_n371_), .ZN(new_n379_));
  NAND3_X1  g242(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g243(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g244(.A(new_n377_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n382_));
  XNOR2_X1  g245(.A(G134gat), .B(G162gat), .ZN(new_n383_));
  XNOR2_X1  g246(.A(new_n383_), .B(G190gat), .ZN(new_n384_));
  INV_X1    g247(.A(new_n384_), .ZN(new_n385_));
  NOR3_X1   g248(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g249(.A1(new_n376_), .A2(new_n379_), .ZN(new_n387_));
  NAND2_X1  g250(.A1(new_n387_), .A2(G218gat), .ZN(new_n388_));
  AOI21_X1  g251(.A(new_n384_), .B1(new_n388_), .B2(new_n380_), .ZN(new_n389_));
  NOR2_X1   g252(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g253(.A(G57gat), .B(G64gat), .ZN(new_n391_));
  INV_X1    g254(.A(G78gat), .ZN(new_n392_));
  NAND3_X1  g255(.A1(new_n391_), .A2(KEYINPUT10), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g256(.A(new_n393_), .B1(new_n392_), .B2(new_n391_), .ZN(new_n394_));
  XNOR2_X1  g257(.A(new_n394_), .B(G71gat), .ZN(new_n395_));
  NAND2_X1  g258(.A1(new_n395_), .A2(KEYINPUT12), .ZN(new_n396_));
  INV_X1    g259(.A(G71gat), .ZN(new_n397_));
  XNOR2_X1  g260(.A(new_n394_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n399_));
  NAND2_X1  g262(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g263(.A1(new_n396_), .A2(new_n400_), .A3(new_n331_), .ZN(new_n401_));
  OAI21_X1  g264(.A(new_n401_), .B1(new_n331_), .B2(new_n398_), .ZN(new_n402_));
  NAND2_X1  g265(.A1(G231gat), .A2(G233gat), .ZN(new_n403_));
  OAI21_X1  g266(.A(new_n402_), .B1(KEYINPUT18), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g267(.A(G127gat), .B(G155gat), .ZN(new_n405_));
  XNOR2_X1  g268(.A(G183gat), .B(G211gat), .ZN(new_n406_));
  XNOR2_X1  g269(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g270(.A1(new_n403_), .A2(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g271(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g272(.A(new_n409_), .B(KEYINPUT19), .Z(new_n410_));
  XNOR2_X1  g273(.A(new_n404_), .B(new_n410_), .ZN(new_n411_));
  NOR2_X1   g274(.A1(new_n390_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g275(.A1(new_n317_), .A2(new_n348_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g276(.A1(new_n413_), .A2(KEYINPUT38), .ZN(new_n414_));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n415_));
  NAND4_X1  g278(.A1(new_n317_), .A2(new_n415_), .A3(new_n348_), .A4(new_n412_), .ZN(new_n416_));
  NAND2_X1  g279(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g280(.A(G1gat), .ZN(new_n418_));
  NAND2_X1  g281(.A1(new_n396_), .A2(new_n400_), .ZN(new_n419_));
  NAND2_X1  g282(.A1(new_n419_), .A2(new_n372_), .ZN(new_n420_));
  INV_X1    g283(.A(new_n366_), .ZN(new_n421_));
  NAND2_X1  g284(.A1(new_n421_), .A2(new_n398_), .ZN(new_n422_));
  OR2_X1    g285(.A1(new_n422_), .A2(KEYINPUT13), .ZN(new_n423_));
  NAND2_X1  g286(.A1(G230gat), .A2(G233gat), .ZN(new_n424_));
  NAND2_X1  g287(.A1(new_n422_), .A2(KEYINPUT13), .ZN(new_n425_));
  NAND4_X1  g288(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  NOR2_X1   g289(.A1(new_n421_), .A2(new_n398_), .ZN(new_n427_));
  INV_X1    g290(.A(new_n422_), .ZN(new_n428_));
  OAI211_X1 g291(.A(G230gat), .B(G233gat), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  AND2_X1   g292(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g293(.A(G176gat), .B(G204gat), .ZN(new_n431_));
  XNOR2_X1  g294(.A(new_n431_), .B(KEYINPUT5), .ZN(new_n432_));
  XNOR2_X1  g295(.A(G120gat), .B(G148gat), .ZN(new_n433_));
  XNOR2_X1  g296(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g297(.A(new_n434_), .B(KEYINPUT6), .ZN(new_n435_));
  OR2_X1    g298(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g299(.A1(new_n426_), .A2(new_n429_), .A3(new_n435_), .ZN(new_n437_));
  NAND2_X1  g300(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g301(.A1(new_n438_), .A2(new_n259_), .ZN(new_n439_));
  NAND3_X1  g302(.A1(new_n417_), .A2(new_n418_), .A3(new_n439_), .ZN(new_n440_));
  NOR3_X1   g303(.A1(new_n413_), .A2(new_n259_), .A3(new_n438_), .ZN(new_n441_));
  OAI21_X1  g304(.A(new_n440_), .B1(new_n418_), .B2(new_n441_), .ZN(G1324gat));
  AND2_X1   g305(.A1(new_n317_), .A2(new_n412_), .ZN(new_n443_));
  INV_X1    g306(.A(new_n438_), .ZN(new_n444_));
  NAND3_X1  g307(.A1(new_n443_), .A2(new_n348_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g308(.A(G8gat), .ZN(new_n446_));
  INV_X1    g309(.A(new_n286_), .ZN(new_n447_));
  NOR3_X1   g310(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g311(.A1(new_n417_), .A2(new_n286_), .A3(new_n444_), .ZN(new_n449_));
  AOI21_X1  g312(.A(new_n448_), .B1(new_n446_), .B2(new_n449_), .ZN(G1325gat));
  INV_X1    g313(.A(new_n192_), .ZN(new_n451_));
  NOR2_X1   g314(.A1(new_n451_), .A2(new_n438_), .ZN(new_n452_));
  AOI21_X1  g315(.A(G15gat), .B1(new_n417_), .B2(new_n452_), .ZN(new_n453_));
  NOR3_X1   g316(.A1(new_n445_), .A2(new_n326_), .A3(new_n314_), .ZN(new_n454_));
  NOR2_X1   g317(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g318(.A(KEYINPUT39), .ZN(new_n456_));
  NAND2_X1  g319(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g320(.A(KEYINPUT39), .B1(new_n453_), .B2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g321(.A1(new_n457_), .A2(new_n458_), .ZN(G1326gat));
  NOR3_X1   g322(.A1(new_n445_), .A2(new_n327_), .A3(new_n239_), .ZN(new_n460_));
  NAND3_X1  g323(.A1(new_n417_), .A2(new_n238_), .A3(new_n444_), .ZN(new_n461_));
  AOI21_X1  g324(.A(new_n460_), .B1(new_n327_), .B2(new_n461_), .ZN(G1327gat));
  NAND2_X1  g325(.A1(new_n310_), .A2(new_n314_), .ZN(new_n463_));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n464_));
  NAND2_X1  g327(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g328(.A1(new_n310_), .A2(new_n314_), .A3(KEYINPUT36), .ZN(new_n466_));
  AOI21_X1  g329(.A(new_n287_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g330(.A(new_n385_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n468_));
  NAND3_X1  g331(.A1(new_n388_), .A2(new_n384_), .A3(new_n380_), .ZN(new_n469_));
  NAND2_X1  g332(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g333(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g334(.A1(new_n471_), .A2(new_n348_), .A3(new_n411_), .ZN(new_n472_));
  XNOR2_X1  g335(.A(new_n472_), .B(KEYINPUT42), .ZN(new_n473_));
  NAND3_X1  g336(.A1(new_n473_), .A2(new_n319_), .A3(new_n439_), .ZN(new_n474_));
  OAI21_X1  g337(.A(KEYINPUT40), .B1(new_n467_), .B2(new_n470_), .ZN(new_n475_));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n476_));
  NAND3_X1  g339(.A1(new_n317_), .A2(new_n476_), .A3(new_n390_), .ZN(new_n477_));
  NAND2_X1  g340(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g341(.A(new_n348_), .ZN(new_n479_));
  NOR2_X1   g342(.A1(new_n438_), .A2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g343(.A1(new_n478_), .A2(new_n411_), .A3(new_n260_), .A4(new_n480_), .ZN(new_n481_));
  AND3_X1   g344(.A1(new_n481_), .A2(KEYINPUT41), .A3(G29gat), .ZN(new_n482_));
  AOI21_X1  g345(.A(KEYINPUT41), .B1(new_n481_), .B2(G29gat), .ZN(new_n483_));
  OAI21_X1  g346(.A(new_n474_), .B1(new_n482_), .B2(new_n483_), .ZN(G1328gat));
  INV_X1    g347(.A(KEYINPUT43), .ZN(new_n485_));
  NAND3_X1  g348(.A1(new_n286_), .A2(new_n485_), .A3(new_n322_), .ZN(new_n486_));
  OAI21_X1  g349(.A(new_n486_), .B1(new_n485_), .B2(new_n322_), .ZN(new_n487_));
  NAND3_X1  g350(.A1(new_n473_), .A2(new_n444_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g351(.A1(new_n478_), .A2(new_n411_), .A3(new_n480_), .ZN(new_n489_));
  OAI21_X1  g352(.A(G36gat), .B1(new_n489_), .B2(new_n447_), .ZN(new_n490_));
  NAND2_X1  g353(.A1(new_n488_), .A2(new_n490_), .ZN(G1329gat));
  INV_X1    g354(.A(G43gat), .ZN(new_n492_));
  NAND3_X1  g355(.A1(new_n473_), .A2(new_n492_), .A3(new_n452_), .ZN(new_n493_));
  OAI21_X1  g356(.A(G43gat), .B1(new_n489_), .B2(new_n314_), .ZN(new_n494_));
  NAND2_X1  g357(.A1(new_n493_), .A2(new_n494_), .ZN(G1330gat));
  OAI21_X1  g358(.A(G50gat), .B1(new_n489_), .B2(new_n239_), .ZN(new_n496_));
  NAND2_X1  g359(.A1(new_n473_), .A2(new_n444_), .ZN(new_n497_));
  OR2_X1    g360(.A1(new_n239_), .A2(G50gat), .ZN(new_n498_));
  OAI21_X1  g361(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(G1331gat));
  NOR2_X1   g362(.A1(new_n444_), .A2(new_n348_), .ZN(new_n500_));
  AND2_X1   g363(.A1(new_n443_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g364(.A1(new_n501_), .A2(new_n260_), .ZN(new_n502_));
  XNOR2_X1  g365(.A(new_n502_), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g366(.A1(new_n501_), .A2(new_n286_), .ZN(new_n504_));
  NAND2_X1  g367(.A1(KEYINPUT44), .A2(G64gat), .ZN(new_n505_));
  NOR2_X1   g368(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g369(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  OR2_X1    g370(.A1(KEYINPUT44), .A2(G64gat), .ZN(new_n508_));
  AOI21_X1  g371(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(G1333gat));
  INV_X1    g372(.A(new_n314_), .ZN(new_n510_));
  AOI21_X1  g373(.A(new_n397_), .B1(new_n501_), .B2(new_n510_), .ZN(new_n511_));
  NAND4_X1  g374(.A1(new_n443_), .A2(KEYINPUT10), .A3(new_n397_), .A4(new_n500_), .ZN(new_n512_));
  OR2_X1    g375(.A1(new_n397_), .A2(KEYINPUT10), .ZN(new_n513_));
  AOI21_X1  g376(.A(new_n451_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g377(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g378(.A1(new_n515_), .A2(KEYINPUT45), .ZN(new_n516_));
  INV_X1    g379(.A(KEYINPUT45), .ZN(new_n517_));
  OAI21_X1  g380(.A(new_n517_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g381(.A1(new_n516_), .A2(new_n518_), .ZN(G1334gat));
  NAND2_X1  g382(.A1(new_n501_), .A2(new_n238_), .ZN(new_n520_));
  XOR2_X1   g383(.A(KEYINPUT46), .B(G78gat), .Z(new_n521_));
  XNOR2_X1  g384(.A(new_n520_), .B(new_n521_), .ZN(G1335gat));
  NAND3_X1  g385(.A1(new_n478_), .A2(new_n411_), .A3(new_n500_), .ZN(new_n523_));
  OAI21_X1  g386(.A(G85gat), .B1(new_n523_), .B2(new_n259_), .ZN(new_n524_));
  INV_X1    g387(.A(new_n411_), .ZN(new_n525_));
  NOR4_X1   g388(.A1(new_n467_), .A2(new_n348_), .A3(new_n470_), .A4(new_n525_), .ZN(new_n526_));
  NAND4_X1  g389(.A1(new_n526_), .A2(new_n254_), .A3(new_n260_), .A4(new_n438_), .ZN(new_n527_));
  NAND2_X1  g390(.A1(new_n524_), .A2(new_n527_), .ZN(G1336gat));
  NOR2_X1   g391(.A1(new_n444_), .A2(new_n447_), .ZN(new_n529_));
  NAND3_X1  g392(.A1(new_n526_), .A2(new_n274_), .A3(new_n529_), .ZN(new_n530_));
  NAND4_X1  g393(.A1(new_n478_), .A2(new_n411_), .A3(new_n286_), .A4(new_n500_), .ZN(new_n531_));
  AND3_X1   g394(.A1(new_n531_), .A2(KEYINPUT47), .A3(G92gat), .ZN(new_n532_));
  AOI21_X1  g395(.A(KEYINPUT47), .B1(new_n531_), .B2(G92gat), .ZN(new_n533_));
  OAI21_X1  g396(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(G1337gat));
  OAI21_X1  g397(.A(G99gat), .B1(new_n523_), .B2(new_n314_), .ZN(new_n535_));
  INV_X1    g398(.A(KEYINPUT48), .ZN(new_n536_));
  NAND2_X1  g399(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g400(.A1(new_n444_), .A2(new_n451_), .ZN(new_n538_));
  NAND3_X1  g401(.A1(new_n526_), .A2(new_n349_), .A3(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g402(.A(new_n539_), .B(KEYINPUT49), .ZN(new_n540_));
  OAI211_X1 g403(.A(KEYINPUT48), .B(G99gat), .C1(new_n523_), .C2(new_n314_), .ZN(new_n541_));
  NAND3_X1  g404(.A1(new_n537_), .A2(new_n540_), .A3(new_n541_), .ZN(G1338gat));
  INV_X1    g405(.A(new_n500_), .ZN(new_n543_));
  AOI211_X1 g406(.A(new_n525_), .B(new_n543_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n544_));
  AOI21_X1  g407(.A(new_n350_), .B1(new_n544_), .B2(new_n238_), .ZN(new_n545_));
  NAND4_X1  g408(.A1(new_n526_), .A2(new_n350_), .A3(new_n238_), .A4(new_n438_), .ZN(new_n546_));
  INV_X1    g409(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g410(.A(KEYINPUT50), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g411(.A(G106gat), .B1(new_n523_), .B2(new_n239_), .ZN(new_n549_));
  INV_X1    g412(.A(KEYINPUT50), .ZN(new_n550_));
  NAND3_X1  g413(.A1(new_n549_), .A2(new_n550_), .A3(new_n546_), .ZN(new_n551_));
  NAND2_X1  g414(.A1(new_n548_), .A2(new_n551_), .ZN(G1339gat));
  INV_X1    g415(.A(KEYINPUT53), .ZN(new_n553_));
  AND3_X1   g416(.A1(new_n420_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n554_));
  OAI21_X1  g417(.A(KEYINPUT52), .B1(new_n554_), .B2(new_n424_), .ZN(new_n555_));
  AOI22_X1  g418(.A1(new_n419_), .A2(new_n372_), .B1(KEYINPUT13), .B2(new_n422_), .ZN(new_n556_));
  AOI21_X1  g419(.A(new_n424_), .B1(new_n556_), .B2(new_n423_), .ZN(new_n557_));
  INV_X1    g420(.A(KEYINPUT52), .ZN(new_n558_));
  NAND2_X1  g421(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g422(.A1(new_n555_), .A2(new_n559_), .A3(new_n426_), .ZN(new_n560_));
  NAND2_X1  g423(.A1(new_n437_), .A2(KEYINPUT51), .ZN(new_n561_));
  INV_X1    g424(.A(KEYINPUT51), .ZN(new_n562_));
  NAND4_X1  g425(.A1(new_n426_), .A2(new_n562_), .A3(new_n429_), .A4(new_n435_), .ZN(new_n563_));
  AOI22_X1  g426(.A1(new_n560_), .A2(new_n434_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g427(.A1(new_n334_), .A2(new_n335_), .ZN(new_n565_));
  AOI21_X1  g428(.A(new_n339_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n566_));
  OAI21_X1  g429(.A(new_n345_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AND2_X1   g430(.A1(new_n567_), .A2(new_n347_), .ZN(new_n568_));
  AOI21_X1  g431(.A(new_n553_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g432(.A(new_n426_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n570_));
  NOR3_X1   g433(.A1(new_n554_), .A2(KEYINPUT52), .A3(new_n424_), .ZN(new_n571_));
  OAI21_X1  g434(.A(new_n434_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g435(.A1(new_n561_), .A2(new_n563_), .ZN(new_n573_));
  AND4_X1   g436(.A1(new_n553_), .A2(new_n572_), .A3(new_n568_), .A4(new_n573_), .ZN(new_n574_));
  OAI21_X1  g437(.A(new_n390_), .B1(new_n569_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g438(.A1(new_n564_), .A2(new_n348_), .ZN(new_n576_));
  NAND2_X1  g439(.A1(new_n438_), .A2(new_n568_), .ZN(new_n577_));
  NAND3_X1  g440(.A1(new_n470_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND3_X1  g441(.A1(new_n575_), .A2(new_n411_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g442(.A1(new_n412_), .A2(new_n479_), .A3(new_n444_), .ZN(new_n580_));
  AOI21_X1  g443(.A(new_n240_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g444(.A1(new_n581_), .A2(new_n260_), .A3(new_n447_), .ZN(new_n582_));
  NOR2_X1   g445(.A1(new_n582_), .A2(new_n479_), .ZN(new_n583_));
  XOR2_X1   g446(.A(KEYINPUT54), .B(G113gat), .Z(new_n584_));
  XNOR2_X1  g447(.A(new_n583_), .B(new_n584_), .ZN(G1340gat));
  NAND2_X1  g448(.A1(KEYINPUT55), .A2(G120gat), .ZN(new_n586_));
  OR3_X1    g449(.A1(new_n582_), .A2(new_n444_), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g450(.A1(KEYINPUT55), .A2(G120gat), .ZN(new_n588_));
  OAI211_X1 g451(.A(new_n586_), .B(new_n588_), .C1(new_n582_), .C2(new_n444_), .ZN(new_n589_));
  AND2_X1   g452(.A1(new_n587_), .A2(new_n589_), .ZN(G1341gat));
  NOR2_X1   g453(.A1(new_n582_), .A2(new_n411_), .ZN(new_n591_));
  XNOR2_X1  g454(.A(new_n591_), .B(new_n138_), .ZN(G1342gat));
  NOR2_X1   g455(.A1(new_n582_), .A2(new_n470_), .ZN(new_n593_));
  XNOR2_X1  g456(.A(new_n593_), .B(new_n140_), .ZN(G1343gat));
  AOI211_X1 g457(.A(new_n239_), .B(new_n510_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n595_));
  NAND3_X1  g458(.A1(new_n595_), .A2(new_n260_), .A3(new_n447_), .ZN(new_n596_));
  NOR2_X1   g459(.A1(new_n596_), .A2(new_n479_), .ZN(new_n597_));
  XNOR2_X1  g460(.A(new_n597_), .B(new_n198_), .ZN(G1344gat));
  NOR2_X1   g461(.A1(new_n596_), .A2(new_n444_), .ZN(new_n599_));
  XNOR2_X1  g462(.A(new_n599_), .B(new_n196_), .ZN(G1345gat));
  NOR2_X1   g463(.A1(new_n596_), .A2(new_n411_), .ZN(new_n601_));
  XNOR2_X1  g464(.A(new_n601_), .B(new_n193_), .ZN(G1346gat));
  NOR2_X1   g465(.A1(new_n596_), .A2(new_n470_), .ZN(new_n603_));
  XNOR2_X1  g466(.A(new_n603_), .B(new_n194_), .ZN(G1347gat));
  NAND3_X1  g467(.A1(new_n581_), .A2(new_n259_), .A3(new_n286_), .ZN(new_n605_));
  NOR2_X1   g468(.A1(new_n605_), .A2(new_n479_), .ZN(new_n606_));
  XNOR2_X1  g469(.A(new_n606_), .B(new_n162_), .ZN(G1348gat));
  INV_X1    g470(.A(KEYINPUT58), .ZN(new_n608_));
  NAND3_X1  g471(.A1(new_n581_), .A2(new_n259_), .A3(new_n529_), .ZN(new_n609_));
  NAND2_X1  g472(.A1(new_n609_), .A2(G176gat), .ZN(new_n610_));
  INV_X1    g473(.A(KEYINPUT56), .ZN(new_n611_));
  NAND2_X1  g474(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g475(.A1(new_n609_), .A2(KEYINPUT56), .A3(G176gat), .ZN(new_n613_));
  NAND2_X1  g476(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g477(.A1(new_n581_), .A2(new_n163_), .A3(new_n259_), .A4(new_n529_), .ZN(new_n615_));
  XNOR2_X1  g478(.A(new_n615_), .B(KEYINPUT57), .ZN(new_n616_));
  OAI21_X1  g479(.A(new_n608_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g480(.A(KEYINPUT57), .ZN(new_n618_));
  XNOR2_X1  g481(.A(new_n615_), .B(new_n618_), .ZN(new_n619_));
  NAND4_X1  g482(.A1(new_n619_), .A2(KEYINPUT58), .A3(new_n612_), .A4(new_n613_), .ZN(new_n620_));
  NAND2_X1  g483(.A1(new_n617_), .A2(new_n620_), .ZN(G1349gat));
  NOR2_X1   g484(.A1(new_n605_), .A2(new_n411_), .ZN(new_n622_));
  XNOR2_X1  g485(.A(new_n622_), .B(new_n174_), .ZN(G1350gat));
  OAI21_X1  g486(.A(G190gat), .B1(new_n605_), .B2(new_n470_), .ZN(new_n624_));
  INV_X1    g487(.A(KEYINPUT59), .ZN(new_n625_));
  OR2_X1    g488(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g489(.A1(new_n605_), .A2(new_n470_), .ZN(new_n627_));
  OAI21_X1  g490(.A(new_n627_), .B1(new_n176_), .B2(new_n175_), .ZN(new_n628_));
  NAND2_X1  g491(.A1(new_n624_), .A2(new_n625_), .ZN(new_n629_));
  NAND3_X1  g492(.A1(new_n626_), .A2(new_n628_), .A3(new_n629_), .ZN(G1351gat));
  NAND2_X1  g493(.A1(new_n579_), .A2(new_n580_), .ZN(new_n631_));
  NAND4_X1  g494(.A1(new_n631_), .A2(new_n259_), .A3(new_n238_), .A4(new_n314_), .ZN(new_n632_));
  OR2_X1    g495(.A1(new_n632_), .A2(KEYINPUT61), .ZN(new_n633_));
  NAND2_X1  g496(.A1(new_n632_), .A2(KEYINPUT61), .ZN(new_n634_));
  AOI21_X1  g497(.A(new_n447_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g498(.A(G197gat), .B1(new_n635_), .B2(new_n348_), .ZN(new_n636_));
  OAI21_X1  g499(.A(KEYINPUT60), .B1(new_n632_), .B2(new_n447_), .ZN(new_n637_));
  INV_X1    g500(.A(KEYINPUT60), .ZN(new_n638_));
  NAND4_X1  g501(.A1(new_n595_), .A2(new_n638_), .A3(new_n259_), .A4(new_n286_), .ZN(new_n639_));
  AND4_X1   g502(.A1(G197gat), .A2(new_n637_), .A3(new_n639_), .A4(new_n348_), .ZN(new_n640_));
  NOR2_X1   g503(.A1(new_n636_), .A2(new_n640_), .ZN(G1352gat));
  AOI21_X1  g504(.A(G204gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n642_));
  NAND2_X1  g505(.A1(new_n642_), .A2(new_n529_), .ZN(new_n643_));
  NAND3_X1  g506(.A1(new_n637_), .A2(new_n639_), .A3(new_n438_), .ZN(new_n644_));
  AND3_X1   g507(.A1(new_n644_), .A2(KEYINPUT62), .A3(G204gat), .ZN(new_n645_));
  AOI21_X1  g508(.A(KEYINPUT62), .B1(new_n644_), .B2(G204gat), .ZN(new_n646_));
  OAI21_X1  g509(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(G1353gat));
  NAND3_X1  g510(.A1(new_n635_), .A2(new_n218_), .A3(new_n525_), .ZN(new_n648_));
  NAND3_X1  g511(.A1(new_n637_), .A2(new_n639_), .A3(new_n525_), .ZN(new_n649_));
  AND3_X1   g512(.A1(new_n649_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n650_));
  AOI21_X1  g513(.A(KEYINPUT63), .B1(new_n649_), .B2(G211gat), .ZN(new_n651_));
  OAI21_X1  g514(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(G1354gat));
  NAND3_X1  g515(.A1(new_n637_), .A2(new_n639_), .A3(new_n390_), .ZN(new_n653_));
  NAND2_X1  g516(.A1(new_n653_), .A2(G218gat), .ZN(new_n654_));
  OAI21_X1  g517(.A(new_n635_), .B1(new_n220_), .B2(new_n219_), .ZN(new_n655_));
  OAI21_X1  g518(.A(new_n654_), .B1(new_n655_), .B2(new_n470_), .ZN(G1355gat));
endmodule


