//Secret key is'1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_c2670" written by ABC on Tue Nov  1 16:41:39 2022

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6,
    G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26,
    G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48,
    G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64,
    G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80,
    G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140,
    G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184,
    G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
    G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210,
    G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245,
    G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
    G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273,
    G274, G275, G276, G277, G278, G279, G452, G483, G543, G559, G567, G651,
    G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966,
    G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078,
    G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435,
    G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3,
    G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24,
    G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44,
    G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62,
    G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78,
    G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94,
    G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138,
    G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196,
    G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208,
    G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243,
    G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255,
    G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271,
    G272, G273, G274, G275, G276, G277, G278, G279, G452, G483, G543, G559,
    G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961,
    G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072,
    G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430,
    G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n383_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n477_, new_n479_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n519_,
    new_n520_, new_n523_, new_n525_, new_n526_, new_n527_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT0), .B(G1083), .ZN(G367));
  XOR2_X1   g005(.A(KEYINPUT1), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  INV_X1    g010(.A(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT3), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(G223));
  NAND3_X1  g021(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n383_));
  XOR2_X1   g022(.A(new_n383_), .B(KEYINPUT4), .Z(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n386_));
  XOR2_X1   g025(.A(new_n386_), .B(KEYINPUT5), .Z(new_n387_));
  INV_X1    g026(.A(new_n387_), .ZN(new_n388_));
  NAND4_X1  g027(.A1(G44), .A2(G82), .A3(G96), .A4(G132), .ZN(new_n389_));
  XNOR2_X1  g028(.A(new_n389_), .B(KEYINPUT6), .ZN(new_n390_));
  INV_X1    g029(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g030(.A1(new_n388_), .A2(new_n391_), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n388_), .A2(G567), .B1(G2106), .B2(new_n391_), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n395_));
  NOR2_X1   g034(.A1(new_n395_), .A2(G2104), .ZN(new_n396_));
  INV_X1    g035(.A(G2104), .ZN(new_n397_));
  NOR2_X1   g036(.A1(new_n397_), .A2(KEYINPUT8), .ZN(new_n398_));
  OAI211_X1 g037(.A(G125), .B(G2105), .C1(new_n396_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g038(.A(KEYINPUT9), .ZN(new_n400_));
  NAND2_X1  g039(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g040(.A1(new_n397_), .A2(KEYINPUT8), .ZN(new_n402_));
  NAND2_X1  g041(.A1(new_n395_), .A2(G2104), .ZN(new_n403_));
  NAND2_X1  g042(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g043(.A1(new_n404_), .A2(KEYINPUT9), .A3(G125), .A4(G2105), .ZN(new_n405_));
  NAND2_X1  g044(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g045(.A1(G113), .A2(G2104), .A3(G2105), .ZN(new_n407_));
  OR2_X1    g046(.A1(KEYINPUT7), .A2(G2105), .ZN(new_n408_));
  NAND2_X1  g047(.A1(KEYINPUT7), .A2(G2105), .ZN(new_n409_));
  AOI22_X1  g048(.A1(new_n402_), .A2(new_n403_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g049(.A(new_n397_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n411_));
  AOI22_X1  g050(.A1(new_n410_), .A2(G137), .B1(new_n411_), .B2(G101), .ZN(new_n412_));
  AND3_X1   g051(.A1(new_n406_), .A2(new_n407_), .A3(new_n412_), .ZN(G160));
  NAND2_X1  g052(.A1(G100), .A2(G2104), .ZN(new_n414_));
  INV_X1    g053(.A(new_n404_), .ZN(new_n415_));
  INV_X1    g054(.A(G136), .ZN(new_n416_));
  OAI21_X1  g055(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g056(.A(KEYINPUT7), .B(G2105), .ZN(new_n418_));
  NAND2_X1  g057(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g058(.A1(G112), .A2(G2104), .ZN(new_n420_));
  INV_X1    g059(.A(G124), .ZN(new_n421_));
  OAI21_X1  g060(.A(new_n420_), .B1(new_n415_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g061(.A1(new_n422_), .A2(G2105), .ZN(new_n423_));
  AND2_X1   g062(.A1(new_n419_), .A2(new_n423_), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT7), .A2(G2105), .ZN(new_n425_));
  NOR2_X1   g064(.A1(KEYINPUT7), .A2(G2105), .ZN(new_n426_));
  OAI211_X1 g065(.A(G102), .B(G2104), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g066(.A1(new_n427_), .A2(KEYINPUT10), .ZN(new_n428_));
  INV_X1    g067(.A(KEYINPUT10), .ZN(new_n429_));
  NAND4_X1  g068(.A1(new_n418_), .A2(new_n429_), .A3(G102), .A4(G2104), .ZN(new_n430_));
  AOI22_X1  g069(.A1(new_n428_), .A2(new_n430_), .B1(new_n410_), .B2(G138), .ZN(new_n431_));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n396_), .C2(new_n398_), .ZN(new_n432_));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n433_));
  NAND2_X1  g072(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g073(.A1(new_n404_), .A2(KEYINPUT11), .A3(G126), .A4(G2105), .ZN(new_n435_));
  NAND2_X1  g074(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g075(.A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n437_));
  NAND3_X1  g076(.A1(new_n431_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g077(.A(new_n438_), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n440_));
  NOR2_X1   g079(.A1(new_n440_), .A2(G75), .ZN(new_n441_));
  NOR2_X1   g080(.A1(G62), .A2(G543), .ZN(new_n442_));
  OAI21_X1  g081(.A(G651), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g082(.A(G651), .ZN(new_n444_));
  NOR2_X1   g083(.A1(new_n440_), .A2(G50), .ZN(new_n445_));
  NOR2_X1   g084(.A1(G88), .A2(G543), .ZN(new_n446_));
  OAI21_X1  g085(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g086(.A1(new_n443_), .A2(new_n447_), .ZN(G166));
  NOR2_X1   g087(.A1(new_n440_), .A2(G76), .ZN(new_n449_));
  NOR2_X1   g088(.A1(G63), .A2(G543), .ZN(new_n450_));
  OAI21_X1  g089(.A(G651), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g090(.A1(new_n440_), .A2(G51), .ZN(new_n452_));
  NOR2_X1   g091(.A1(G89), .A2(G543), .ZN(new_n453_));
  OAI21_X1  g092(.A(new_n444_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g093(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g094(.A1(new_n455_), .A2(KEYINPUT12), .ZN(new_n456_));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n457_));
  NAND3_X1  g096(.A1(new_n451_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g097(.A1(new_n456_), .A2(new_n458_), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  NAND3_X1  g099(.A1(new_n440_), .A2(G64), .A3(G651), .ZN(new_n461_));
  XOR2_X1   g100(.A(new_n461_), .B(KEYINPUT13), .Z(new_n462_));
  MUX2_X1   g101(.A(G90), .B(G52), .S(G543), .Z(new_n463_));
  AOI21_X1  g102(.A(new_n462_), .B1(new_n444_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g103(.A1(G77), .A2(G543), .A3(G651), .ZN(new_n465_));
  XOR2_X1   g104(.A(new_n465_), .B(KEYINPUT14), .Z(new_n466_));
  NAND2_X1  g105(.A1(new_n464_), .A2(new_n466_), .ZN(G301));
  XOR2_X1   g106(.A(G301), .B(KEYINPUT15), .Z(G171));
  NAND3_X1  g107(.A1(new_n444_), .A2(G43), .A3(G543), .ZN(new_n469_));
  XOR2_X1   g108(.A(new_n469_), .B(KEYINPUT16), .Z(new_n470_));
  AND3_X1   g109(.A1(G68), .A2(G543), .A3(G651), .ZN(new_n471_));
  MUX2_X1   g110(.A(G81), .B(G56), .S(G651), .Z(new_n472_));
  AOI21_X1  g111(.A(new_n471_), .B1(new_n472_), .B2(new_n440_), .ZN(new_n473_));
  NAND2_X1  g112(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g113(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g114(.A1(new_n475_), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n477_));
  NAND2_X1  g116(.A1(new_n477_), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n479_));
  NAND2_X1  g118(.A1(new_n477_), .A2(new_n479_), .ZN(G188));
  NOR2_X1   g119(.A1(new_n440_), .A2(G78), .ZN(new_n481_));
  NOR2_X1   g120(.A1(G65), .A2(G543), .ZN(new_n482_));
  OAI21_X1  g121(.A(G651), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g122(.A1(new_n440_), .A2(G53), .ZN(new_n484_));
  NOR2_X1   g123(.A1(G91), .A2(G543), .ZN(new_n485_));
  OAI21_X1  g124(.A(new_n444_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g125(.A1(new_n483_), .A2(new_n486_), .ZN(G299));
  INV_X1    g126(.A(G166), .ZN(G303));
  NOR2_X1   g127(.A1(new_n444_), .A2(G74), .ZN(new_n489_));
  NOR2_X1   g128(.A1(G49), .A2(G651), .ZN(new_n490_));
  OAI21_X1  g129(.A(G543), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g130(.A(new_n491_), .ZN(new_n492_));
  NOR3_X1   g131(.A1(G87), .A2(G543), .A3(G651), .ZN(new_n493_));
  NOR2_X1   g132(.A1(new_n492_), .A2(new_n493_), .ZN(G288));
  AND3_X1   g133(.A1(new_n440_), .A2(G61), .A3(G651), .ZN(new_n495_));
  MUX2_X1   g134(.A(G86), .B(G48), .S(G543), .Z(new_n496_));
  AOI21_X1  g135(.A(new_n495_), .B1(new_n496_), .B2(new_n444_), .ZN(new_n497_));
  NAND3_X1  g136(.A1(G73), .A2(G543), .A3(G651), .ZN(new_n498_));
  XNOR2_X1  g137(.A(new_n498_), .B(KEYINPUT17), .ZN(new_n499_));
  NAND2_X1  g138(.A1(new_n497_), .A2(new_n499_), .ZN(G305));
  NOR2_X1   g139(.A1(new_n440_), .A2(G72), .ZN(new_n501_));
  NOR2_X1   g140(.A1(G60), .A2(G543), .ZN(new_n502_));
  OAI21_X1  g141(.A(G651), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g142(.A1(new_n440_), .A2(G47), .ZN(new_n504_));
  NOR2_X1   g143(.A1(G85), .A2(G543), .ZN(new_n505_));
  OAI21_X1  g144(.A(new_n444_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AND2_X1   g145(.A1(new_n503_), .A2(new_n506_), .ZN(G290));
  NAND2_X1  g146(.A1(G301), .A2(G868), .ZN(new_n508_));
  AND3_X1   g147(.A1(G79), .A2(G543), .A3(G651), .ZN(new_n509_));
  NAND2_X1  g148(.A1(G66), .A2(G651), .ZN(new_n510_));
  INV_X1    g149(.A(G92), .ZN(new_n511_));
  OAI21_X1  g150(.A(new_n510_), .B1(new_n511_), .B2(G651), .ZN(new_n512_));
  AOI21_X1  g151(.A(new_n509_), .B1(new_n512_), .B2(new_n440_), .ZN(new_n513_));
  XOR2_X1   g152(.A(new_n513_), .B(KEYINPUT18), .Z(new_n514_));
  NAND3_X1  g153(.A1(new_n444_), .A2(G54), .A3(G543), .ZN(new_n515_));
  AND2_X1   g154(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g155(.A(new_n508_), .B1(new_n516_), .B2(G868), .ZN(G284));
  OAI21_X1  g156(.A(new_n508_), .B1(new_n516_), .B2(G868), .ZN(G321));
  INV_X1    g157(.A(G868), .ZN(new_n519_));
  NAND2_X1  g158(.A1(G299), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g159(.A(new_n520_), .B1(G168), .B2(new_n519_), .ZN(G297));
  OAI21_X1  g160(.A(new_n520_), .B1(G168), .B2(new_n519_), .ZN(G280));
  INV_X1    g161(.A(G559), .ZN(new_n523_));
  OAI21_X1  g162(.A(new_n516_), .B1(new_n523_), .B2(G860), .ZN(G148));
  NAND2_X1  g163(.A1(new_n474_), .A2(new_n519_), .ZN(new_n525_));
  NAND2_X1  g164(.A1(new_n514_), .A2(new_n515_), .ZN(new_n526_));
  NOR2_X1   g165(.A1(new_n526_), .A2(G559), .ZN(new_n527_));
  OAI21_X1  g166(.A(new_n525_), .B1(new_n527_), .B2(new_n519_), .ZN(G282));
  OAI21_X1  g167(.A(new_n525_), .B1(new_n527_), .B2(new_n519_), .ZN(G323));
  INV_X1    g168(.A(KEYINPUT19), .ZN(new_n530_));
  NAND2_X1  g169(.A1(new_n404_), .A2(new_n418_), .ZN(new_n531_));
  INV_X1    g170(.A(G135), .ZN(new_n532_));
  OAI21_X1  g171(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g172(.A1(new_n410_), .A2(KEYINPUT19), .A3(G135), .ZN(new_n534_));
  NAND2_X1  g173(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g174(.A1(new_n404_), .A2(G123), .A3(G2105), .ZN(new_n536_));
  NAND2_X1  g175(.A1(new_n411_), .A2(G99), .ZN(new_n537_));
  NAND3_X1  g176(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g177(.A1(G111), .A2(G2104), .A3(G2105), .ZN(new_n539_));
  INV_X1    g178(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g179(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g180(.A(new_n541_), .ZN(new_n542_));
  OR2_X1    g181(.A1(new_n542_), .A2(G2096), .ZN(new_n543_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n544_));
  OR3_X1    g183(.A1(new_n404_), .A2(new_n544_), .A3(G2105), .ZN(new_n545_));
  OAI21_X1  g184(.A(new_n544_), .B1(new_n404_), .B2(G2105), .ZN(new_n546_));
  NAND3_X1  g185(.A1(new_n545_), .A2(new_n411_), .A3(new_n546_), .ZN(new_n547_));
  XOR2_X1   g186(.A(new_n547_), .B(G2100), .Z(new_n548_));
  NAND2_X1  g187(.A1(new_n542_), .A2(G2096), .ZN(new_n549_));
  NAND3_X1  g188(.A1(new_n543_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  XOR2_X1   g189(.A(new_n550_), .B(KEYINPUT21), .Z(G156));
  XNOR2_X1  g190(.A(G2427), .B(G2430), .ZN(new_n552_));
  XNOR2_X1  g191(.A(new_n552_), .B(KEYINPUT23), .ZN(new_n553_));
  INV_X1    g192(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g193(.A(G2435), .B(G2438), .Z(new_n555_));
  OR2_X1    g194(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g195(.A1(new_n554_), .A2(new_n555_), .ZN(new_n557_));
  NAND3_X1  g196(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT22), .ZN(new_n558_));
  XOR2_X1   g197(.A(G2443), .B(G2446), .Z(new_n559_));
  XNOR2_X1  g198(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n561_));
  XNOR2_X1  g200(.A(new_n561_), .B(KEYINPUT24), .ZN(new_n562_));
  XOR2_X1   g201(.A(G1341), .B(G1348), .Z(new_n563_));
  XNOR2_X1  g202(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g203(.A(new_n560_), .B(new_n564_), .ZN(new_n565_));
  AND2_X1   g204(.A1(new_n565_), .A2(G14), .ZN(G401));
  XOR2_X1   g205(.A(G2067), .B(G2678), .Z(new_n567_));
  XNOR2_X1  g206(.A(new_n567_), .B(KEYINPUT25), .ZN(new_n568_));
  XNOR2_X1  g207(.A(G2072), .B(G2078), .ZN(new_n569_));
  XNOR2_X1  g208(.A(G2084), .B(G2090), .ZN(new_n570_));
  XNOR2_X1  g209(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g210(.A(new_n568_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g211(.A(G2096), .B(G2100), .Z(new_n573_));
  XNOR2_X1  g212(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g213(.A(new_n574_), .B(KEYINPUT26), .ZN(G227));
  XOR2_X1   g214(.A(G1961), .B(G1966), .Z(new_n576_));
  XOR2_X1   g215(.A(new_n576_), .B(KEYINPUT27), .Z(new_n577_));
  XNOR2_X1  g216(.A(G1971), .B(G1976), .ZN(new_n578_));
  XOR2_X1   g217(.A(G1956), .B(G2474), .Z(new_n579_));
  INV_X1    g218(.A(new_n579_), .ZN(new_n580_));
  NOR3_X1   g219(.A1(new_n577_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  OAI21_X1  g220(.A(new_n580_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n582_));
  NAND2_X1  g221(.A1(new_n576_), .A2(new_n578_), .ZN(new_n583_));
  AOI21_X1  g222(.A(KEYINPUT27), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  OAI22_X1  g223(.A1(new_n581_), .A2(new_n584_), .B1(new_n583_), .B2(new_n579_), .ZN(new_n585_));
  XNOR2_X1  g224(.A(G1991), .B(G1996), .ZN(new_n586_));
  XNOR2_X1  g225(.A(new_n586_), .B(KEYINPUT28), .ZN(new_n587_));
  XOR2_X1   g226(.A(G1981), .B(G1986), .Z(new_n588_));
  XNOR2_X1  g227(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g228(.A(new_n585_), .B(new_n589_), .ZN(G229));
  NAND3_X1  g229(.A1(G116), .A2(G2104), .A3(G2105), .ZN(new_n591_));
  XOR2_X1   g230(.A(new_n591_), .B(KEYINPUT32), .Z(new_n592_));
  NAND2_X1  g231(.A1(new_n411_), .A2(G104), .ZN(new_n593_));
  AOI22_X1  g232(.A1(new_n418_), .A2(G140), .B1(G128), .B2(G2105), .ZN(new_n594_));
  OAI211_X1 g233(.A(new_n592_), .B(new_n593_), .C1(new_n594_), .C2(new_n415_), .ZN(new_n595_));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n596_));
  NAND2_X1  g235(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g236(.A1(G128), .A2(G2105), .ZN(new_n598_));
  NOR2_X1   g237(.A1(new_n425_), .A2(new_n426_), .ZN(new_n599_));
  INV_X1    g238(.A(G140), .ZN(new_n600_));
  OAI21_X1  g239(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g240(.A1(new_n601_), .A2(new_n404_), .ZN(new_n602_));
  NAND4_X1  g241(.A1(new_n602_), .A2(KEYINPUT33), .A3(new_n592_), .A4(new_n593_), .ZN(new_n603_));
  NAND2_X1  g242(.A1(new_n597_), .A2(new_n603_), .ZN(new_n604_));
  MUX2_X1   g243(.A(G26), .B(new_n604_), .S(G29), .Z(new_n605_));
  XNOR2_X1  g244(.A(new_n605_), .B(G2067), .ZN(new_n606_));
  INV_X1    g245(.A(G16), .ZN(new_n607_));
  NAND2_X1  g246(.A1(new_n607_), .A2(G21), .ZN(new_n608_));
  OAI21_X1  g247(.A(new_n608_), .B1(G168), .B2(new_n607_), .ZN(new_n609_));
  XNOR2_X1  g248(.A(new_n609_), .B(G1966), .ZN(new_n610_));
  NOR2_X1   g249(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g250(.A(G29), .ZN(new_n612_));
  NAND2_X1  g251(.A1(new_n612_), .A2(G27), .ZN(new_n613_));
  OAI21_X1  g252(.A(new_n613_), .B1(G164), .B2(new_n612_), .ZN(new_n614_));
  XNOR2_X1  g253(.A(new_n614_), .B(G2078), .ZN(new_n615_));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n616_));
  NAND2_X1  g255(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g256(.A(G2078), .ZN(new_n618_));
  XNOR2_X1  g257(.A(new_n614_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g258(.A1(new_n619_), .A2(KEYINPUT34), .ZN(new_n620_));
  NAND2_X1  g259(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g260(.A1(new_n607_), .A2(G4), .ZN(new_n622_));
  AOI21_X1  g261(.A(new_n622_), .B1(new_n526_), .B2(G16), .ZN(new_n623_));
  INV_X1    g262(.A(G1348), .ZN(new_n624_));
  XNOR2_X1  g263(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NAND2_X1  g264(.A1(new_n607_), .A2(G20), .ZN(new_n626_));
  INV_X1    g265(.A(G299), .ZN(new_n627_));
  OAI21_X1  g266(.A(new_n626_), .B1(new_n627_), .B2(new_n607_), .ZN(new_n628_));
  XNOR2_X1  g267(.A(new_n628_), .B(G1956), .ZN(new_n629_));
  NAND2_X1  g268(.A1(new_n607_), .A2(G19), .ZN(new_n630_));
  OAI21_X1  g269(.A(new_n630_), .B1(new_n475_), .B2(new_n607_), .ZN(new_n631_));
  XNOR2_X1  g270(.A(new_n631_), .B(G1341), .ZN(new_n632_));
  NOR3_X1   g271(.A1(new_n625_), .A2(new_n629_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g272(.A1(new_n607_), .A2(G5), .ZN(new_n634_));
  INV_X1    g273(.A(G301), .ZN(new_n635_));
  OAI21_X1  g274(.A(new_n634_), .B1(new_n635_), .B2(new_n607_), .ZN(new_n636_));
  INV_X1    g275(.A(G1961), .ZN(new_n637_));
  XNOR2_X1  g276(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND4_X1  g277(.A1(new_n611_), .A2(new_n621_), .A3(new_n633_), .A4(new_n638_), .ZN(new_n639_));
  NAND2_X1  g278(.A1(new_n419_), .A2(new_n423_), .ZN(new_n640_));
  NAND2_X1  g279(.A1(new_n640_), .A2(G29), .ZN(new_n641_));
  NAND2_X1  g280(.A1(new_n612_), .A2(G35), .ZN(new_n642_));
  AND2_X1   g281(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g282(.A(G2090), .ZN(new_n644_));
  NOR2_X1   g283(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g284(.A1(new_n612_), .A2(G32), .ZN(new_n646_));
  AOI22_X1  g285(.A1(new_n418_), .A2(G141), .B1(G129), .B2(G2105), .ZN(new_n647_));
  NOR2_X1   g286(.A1(new_n647_), .A2(new_n415_), .ZN(new_n648_));
  NAND2_X1  g287(.A1(new_n411_), .A2(G105), .ZN(new_n649_));
  INV_X1    g288(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n651_));
  XOR2_X1   g290(.A(new_n651_), .B(KEYINPUT31), .Z(new_n652_));
  NOR3_X1   g291(.A1(new_n648_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g292(.A(new_n646_), .B1(new_n653_), .B2(new_n612_), .ZN(new_n654_));
  INV_X1    g293(.A(G1996), .ZN(new_n655_));
  XNOR2_X1  g294(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g295(.A(new_n643_), .ZN(new_n657_));
  OAI21_X1  g296(.A(new_n656_), .B1(G2090), .B2(new_n657_), .ZN(new_n658_));
  NOR3_X1   g297(.A1(new_n639_), .A2(new_n645_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g298(.A1(new_n612_), .A2(G25), .ZN(new_n660_));
  AOI22_X1  g299(.A1(new_n418_), .A2(G131), .B1(G119), .B2(G2105), .ZN(new_n661_));
  NOR2_X1   g300(.A1(new_n661_), .A2(new_n415_), .ZN(new_n662_));
  AOI22_X1  g301(.A1(new_n418_), .A2(G95), .B1(G107), .B2(G2105), .ZN(new_n663_));
  NOR2_X1   g302(.A1(new_n663_), .A2(new_n397_), .ZN(new_n664_));
  NOR2_X1   g303(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g304(.A(new_n660_), .B1(new_n665_), .B2(new_n612_), .ZN(new_n666_));
  XNOR2_X1  g305(.A(KEYINPUT38), .B(G1991), .ZN(new_n667_));
  XNOR2_X1  g306(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  NAND2_X1  g307(.A1(new_n607_), .A2(G6), .ZN(new_n669_));
  INV_X1    g308(.A(G305), .ZN(new_n670_));
  OAI21_X1  g309(.A(new_n669_), .B1(new_n670_), .B2(new_n607_), .ZN(new_n671_));
  INV_X1    g310(.A(G1981), .ZN(new_n672_));
  XNOR2_X1  g311(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  MUX2_X1   g312(.A(G24), .B(G290), .S(G16), .Z(new_n674_));
  NAND2_X1  g313(.A1(new_n674_), .A2(G1986), .ZN(new_n675_));
  NAND3_X1  g314(.A1(new_n668_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g315(.A(KEYINPUT36), .B(G23), .ZN(new_n677_));
  NOR2_X1   g316(.A1(new_n677_), .A2(G16), .ZN(new_n678_));
  XNOR2_X1  g317(.A(new_n678_), .B(KEYINPUT37), .ZN(new_n679_));
  AOI21_X1  g318(.A(new_n679_), .B1(G16), .B2(G288), .ZN(new_n680_));
  XNOR2_X1  g319(.A(new_n680_), .B(G1976), .ZN(new_n681_));
  OAI21_X1  g320(.A(new_n681_), .B1(G1986), .B2(new_n674_), .ZN(new_n682_));
  NAND2_X1  g321(.A1(new_n607_), .A2(G22), .ZN(new_n683_));
  OAI21_X1  g322(.A(new_n683_), .B1(G166), .B2(new_n607_), .ZN(new_n684_));
  XNOR2_X1  g323(.A(new_n684_), .B(G1971), .ZN(new_n685_));
  NOR3_X1   g324(.A1(new_n676_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n687_));
  OR2_X1    g326(.A1(new_n687_), .A2(G34), .ZN(new_n688_));
  NAND2_X1  g327(.A1(new_n687_), .A2(G34), .ZN(new_n689_));
  AOI21_X1  g328(.A(G29), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g329(.A1(new_n406_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n691_));
  AOI21_X1  g330(.A(new_n690_), .B1(new_n691_), .B2(G29), .ZN(new_n692_));
  XNOR2_X1  g331(.A(new_n692_), .B(G2084), .ZN(new_n693_));
  NAND2_X1  g332(.A1(new_n541_), .A2(G29), .ZN(new_n694_));
  OAI21_X1  g333(.A(new_n694_), .B1(G28), .B2(G29), .ZN(new_n695_));
  NAND2_X1  g334(.A1(new_n612_), .A2(G33), .ZN(new_n696_));
  XNOR2_X1  g335(.A(new_n696_), .B(KEYINPUT30), .ZN(new_n697_));
  AOI22_X1  g336(.A1(new_n418_), .A2(G103), .B1(G115), .B2(G2105), .ZN(new_n698_));
  AOI22_X1  g337(.A1(new_n418_), .A2(G139), .B1(G127), .B2(G2105), .ZN(new_n699_));
  OAI22_X1  g338(.A1(new_n397_), .A2(new_n698_), .B1(new_n699_), .B2(new_n415_), .ZN(new_n700_));
  INV_X1    g339(.A(new_n700_), .ZN(new_n701_));
  OAI21_X1  g340(.A(new_n697_), .B1(new_n701_), .B2(new_n612_), .ZN(new_n702_));
  XNOR2_X1  g341(.A(new_n702_), .B(G2072), .ZN(new_n703_));
  NAND3_X1  g342(.A1(KEYINPUT35), .A2(G11), .A3(G868), .ZN(new_n704_));
  OAI21_X1  g343(.A(new_n704_), .B1(KEYINPUT35), .B2(G11), .ZN(new_n705_));
  NOR3_X1   g344(.A1(new_n695_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  NAND4_X1  g345(.A1(new_n659_), .A2(new_n686_), .A3(new_n693_), .A4(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g346(.A(new_n707_), .B(KEYINPUT39), .ZN(G311));
  INV_X1    g347(.A(KEYINPUT39), .ZN(new_n709_));
  XNOR2_X1  g348(.A(new_n707_), .B(new_n709_), .ZN(G150));
  AOI21_X1  g349(.A(new_n475_), .B1(new_n516_), .B2(G559), .ZN(new_n711_));
  NOR3_X1   g350(.A1(new_n526_), .A2(new_n523_), .A3(new_n474_), .ZN(new_n712_));
  NOR3_X1   g351(.A1(new_n711_), .A2(new_n712_), .A3(G860), .ZN(new_n713_));
  MUX2_X1   g352(.A(G93), .B(G55), .S(G543), .Z(new_n714_));
  NAND2_X1  g353(.A1(new_n714_), .A2(new_n444_), .ZN(new_n715_));
  AND2_X1   g354(.A1(G80), .A2(G543), .ZN(new_n716_));
  AOI21_X1  g355(.A(new_n716_), .B1(G67), .B2(new_n440_), .ZN(new_n717_));
  OAI211_X1 g356(.A(new_n715_), .B(KEYINPUT40), .C1(new_n717_), .C2(new_n444_), .ZN(new_n718_));
  INV_X1    g357(.A(KEYINPUT40), .ZN(new_n719_));
  NAND4_X1  g358(.A1(new_n719_), .A2(new_n444_), .A3(G55), .A4(G543), .ZN(new_n720_));
  NAND2_X1  g359(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g360(.A(new_n713_), .B(new_n721_), .ZN(G145));
  XNOR2_X1  g361(.A(KEYINPUT44), .B(G37), .ZN(new_n723_));
  OAI21_X1  g362(.A(new_n547_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n724_));
  INV_X1    g363(.A(new_n547_), .ZN(new_n725_));
  AOI22_X1  g364(.A1(new_n533_), .A2(new_n534_), .B1(G99), .B2(new_n411_), .ZN(new_n726_));
  NAND4_X1  g365(.A1(new_n725_), .A2(new_n726_), .A3(new_n539_), .A4(new_n536_), .ZN(new_n727_));
  NAND2_X1  g366(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g367(.A1(G160), .A2(new_n640_), .ZN(new_n729_));
  NAND2_X1  g368(.A1(G162), .A2(new_n691_), .ZN(new_n730_));
  NAND2_X1  g369(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g370(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g371(.A(KEYINPUT43), .ZN(new_n733_));
  NAND4_X1  g372(.A1(new_n724_), .A2(new_n729_), .A3(new_n730_), .A4(new_n727_), .ZN(new_n734_));
  AND3_X1   g373(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g374(.A(new_n733_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n736_));
  NOR2_X1   g375(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g376(.A1(new_n701_), .A2(new_n437_), .A3(new_n436_), .A4(new_n431_), .ZN(new_n738_));
  NAND2_X1  g377(.A1(new_n438_), .A2(new_n700_), .ZN(new_n739_));
  AOI21_X1  g378(.A(KEYINPUT41), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g379(.A(new_n740_), .ZN(new_n741_));
  NAND3_X1  g380(.A1(new_n653_), .A2(new_n597_), .A3(new_n603_), .ZN(new_n742_));
  INV_X1    g381(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g382(.A(new_n653_), .B1(new_n597_), .B2(new_n603_), .ZN(new_n744_));
  NOR2_X1   g383(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g384(.A1(new_n738_), .A2(new_n739_), .A3(KEYINPUT41), .ZN(new_n746_));
  NAND3_X1  g385(.A1(new_n741_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g386(.A(new_n653_), .ZN(new_n748_));
  NAND2_X1  g387(.A1(new_n604_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g388(.A1(new_n749_), .A2(new_n742_), .ZN(new_n750_));
  AND3_X1   g389(.A1(new_n738_), .A2(KEYINPUT41), .A3(new_n739_), .ZN(new_n751_));
  OAI21_X1  g390(.A(new_n750_), .B1(new_n751_), .B2(new_n740_), .ZN(new_n752_));
  NAND3_X1  g391(.A1(new_n404_), .A2(G130), .A3(G2105), .ZN(new_n753_));
  XOR2_X1   g392(.A(new_n753_), .B(KEYINPUT42), .Z(new_n754_));
  NAND3_X1  g393(.A1(G118), .A2(G2104), .A3(G2105), .ZN(new_n755_));
  AOI22_X1  g394(.A1(new_n410_), .A2(G142), .B1(new_n411_), .B2(G106), .ZN(new_n756_));
  NAND3_X1  g395(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g396(.A(new_n757_), .B(new_n665_), .ZN(new_n758_));
  AND3_X1   g397(.A1(new_n747_), .A2(new_n752_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g398(.A(new_n758_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n760_));
  OAI21_X1  g399(.A(new_n737_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g400(.A1(new_n747_), .A2(new_n752_), .ZN(new_n762_));
  INV_X1    g401(.A(new_n758_), .ZN(new_n763_));
  NAND2_X1  g402(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g403(.A(new_n734_), .ZN(new_n765_));
  AOI22_X1  g404(.A1(new_n724_), .A2(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n766_));
  OAI21_X1  g405(.A(KEYINPUT43), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g406(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n768_));
  NAND2_X1  g407(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g408(.A1(new_n747_), .A2(new_n752_), .A3(new_n758_), .ZN(new_n770_));
  NAND3_X1  g409(.A1(new_n764_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g410(.A(new_n723_), .B1(new_n761_), .B2(new_n771_), .ZN(G395));
  XNOR2_X1  g411(.A(new_n526_), .B(G299), .ZN(new_n773_));
  XNOR2_X1  g412(.A(new_n721_), .B(new_n474_), .ZN(new_n774_));
  XNOR2_X1  g413(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  NAND2_X1  g414(.A1(new_n775_), .A2(KEYINPUT45), .ZN(new_n776_));
  INV_X1    g415(.A(new_n527_), .ZN(new_n777_));
  NAND2_X1  g416(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g417(.A1(new_n775_), .A2(KEYINPUT45), .A3(new_n527_), .ZN(new_n779_));
  INV_X1    g418(.A(KEYINPUT45), .ZN(new_n780_));
  OAI21_X1  g419(.A(new_n780_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n781_));
  NAND3_X1  g420(.A1(new_n778_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g421(.A(G305), .B(G290), .ZN(new_n783_));
  XNOR2_X1  g422(.A(G288), .B(G166), .ZN(new_n784_));
  XNOR2_X1  g423(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  NAND2_X1  g424(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g425(.A(new_n785_), .ZN(new_n787_));
  NAND4_X1  g426(.A1(new_n778_), .A2(new_n787_), .A3(new_n779_), .A4(new_n781_), .ZN(new_n788_));
  NAND3_X1  g427(.A1(new_n786_), .A2(G868), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g428(.A1(new_n718_), .A2(new_n519_), .A3(new_n720_), .ZN(new_n790_));
  NAND2_X1  g429(.A1(new_n789_), .A2(new_n790_), .ZN(G331));
  NAND2_X1  g430(.A1(G331), .A2(KEYINPUT46), .ZN(new_n792_));
  INV_X1    g431(.A(KEYINPUT46), .ZN(new_n793_));
  NAND3_X1  g432(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g433(.A1(new_n792_), .A2(new_n794_), .ZN(G295));
  XNOR2_X1  g434(.A(G301), .B(G286), .ZN(new_n796_));
  XNOR2_X1  g435(.A(new_n775_), .B(new_n796_), .ZN(new_n797_));
  OR2_X1    g436(.A1(new_n797_), .A2(new_n787_), .ZN(new_n798_));
  INV_X1    g437(.A(new_n723_), .ZN(new_n799_));
  NAND2_X1  g438(.A1(new_n797_), .A2(new_n787_), .ZN(new_n800_));
  NAND3_X1  g439(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g440(.A(new_n801_), .ZN(G397));
  INV_X1    g441(.A(KEYINPUT57), .ZN(new_n803_));
  INV_X1    g442(.A(KEYINPUT56), .ZN(new_n804_));
  INV_X1    g443(.A(G1384), .ZN(new_n805_));
  NAND2_X1  g444(.A1(new_n438_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g445(.A1(new_n406_), .A2(G40), .A3(new_n407_), .A4(new_n412_), .ZN(new_n807_));
  OAI21_X1  g446(.A(new_n624_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g447(.A(new_n807_), .ZN(new_n809_));
  INV_X1    g448(.A(G2067), .ZN(new_n810_));
  NAND4_X1  g449(.A1(new_n809_), .A2(new_n805_), .A3(new_n810_), .A4(new_n438_), .ZN(new_n811_));
  NAND2_X1  g450(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g451(.A(new_n804_), .B1(new_n812_), .B2(new_n516_), .ZN(new_n813_));
  AOI211_X1 g452(.A(KEYINPUT56), .B(new_n526_), .C1(new_n808_), .C2(new_n811_), .ZN(new_n814_));
  NOR2_X1   g453(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g454(.A1(G160), .A2(G40), .A3(new_n805_), .A4(new_n438_), .ZN(new_n816_));
  INV_X1    g455(.A(G1956), .ZN(new_n817_));
  NAND2_X1  g456(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AND2_X1   g457(.A1(new_n438_), .A2(new_n805_), .ZN(new_n819_));
  INV_X1    g458(.A(G2072), .ZN(new_n820_));
  NAND3_X1  g459(.A1(new_n819_), .A2(new_n820_), .A3(new_n809_), .ZN(new_n821_));
  NAND2_X1  g460(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g461(.A1(new_n822_), .A2(new_n627_), .ZN(new_n823_));
  NAND3_X1  g462(.A1(new_n818_), .A2(new_n821_), .A3(G299), .ZN(new_n824_));
  NAND2_X1  g463(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g464(.A(new_n803_), .B1(new_n815_), .B2(new_n825_), .ZN(new_n826_));
  AND3_X1   g465(.A1(new_n818_), .A2(new_n821_), .A3(G299), .ZN(new_n827_));
  AOI21_X1  g466(.A(G299), .B1(new_n818_), .B2(new_n821_), .ZN(new_n828_));
  NOR2_X1   g467(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g468(.A(new_n829_), .B(KEYINPUT57), .C1(new_n813_), .C2(new_n814_), .ZN(new_n830_));
  NAND2_X1  g469(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g470(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g471(.A1(new_n812_), .A2(new_n516_), .ZN(new_n833_));
  NAND3_X1  g472(.A1(new_n808_), .A2(new_n811_), .A3(new_n526_), .ZN(new_n834_));
  NAND3_X1  g473(.A1(new_n833_), .A2(new_n475_), .A3(new_n834_), .ZN(new_n835_));
  XOR2_X1   g474(.A(KEYINPUT59), .B(G1341), .Z(new_n836_));
  NAND2_X1  g475(.A1(new_n816_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g476(.A(KEYINPUT60), .ZN(new_n838_));
  NAND2_X1  g477(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g478(.A1(new_n816_), .A2(KEYINPUT60), .A3(new_n836_), .ZN(new_n840_));
  NOR2_X1   g479(.A1(new_n806_), .A2(new_n807_), .ZN(new_n841_));
  AOI22_X1  g480(.A1(new_n839_), .A2(new_n840_), .B1(new_n655_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g481(.A(new_n823_), .B1(new_n835_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g482(.A(new_n832_), .B1(new_n843_), .B2(new_n824_), .ZN(new_n844_));
  NOR2_X1   g483(.A1(new_n823_), .A2(KEYINPUT58), .ZN(new_n845_));
  OAI21_X1  g484(.A(new_n831_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g485(.A(G1976), .B1(new_n492_), .B2(new_n493_), .ZN(new_n847_));
  OAI211_X1 g486(.A(G8), .B(new_n847_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n848_));
  NAND2_X1  g487(.A1(new_n848_), .A2(KEYINPUT53), .ZN(new_n849_));
  INV_X1    g488(.A(G1976), .ZN(new_n850_));
  NAND4_X1  g489(.A1(new_n816_), .A2(G8), .A3(new_n850_), .A4(G288), .ZN(new_n851_));
  INV_X1    g490(.A(KEYINPUT53), .ZN(new_n852_));
  NAND4_X1  g491(.A1(new_n816_), .A2(new_n852_), .A3(G8), .A4(new_n847_), .ZN(new_n853_));
  NAND3_X1  g492(.A1(new_n849_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g493(.A(G8), .ZN(new_n855_));
  NOR2_X1   g494(.A1(new_n841_), .A2(new_n855_), .ZN(new_n856_));
  XOR2_X1   g495(.A(KEYINPUT51), .B(G1981), .Z(new_n857_));
  XNOR2_X1  g496(.A(G305), .B(new_n857_), .ZN(new_n858_));
  NAND2_X1  g497(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g498(.A(KEYINPUT52), .ZN(new_n860_));
  AOI21_X1  g499(.A(new_n860_), .B1(G286), .B2(G8), .ZN(new_n861_));
  AOI211_X1 g500(.A(KEYINPUT52), .B(new_n855_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n862_));
  NOR2_X1   g501(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g502(.A(G1966), .ZN(new_n864_));
  OAI21_X1  g503(.A(new_n864_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n865_));
  INV_X1    g504(.A(G2084), .ZN(new_n866_));
  NAND4_X1  g505(.A1(new_n809_), .A2(new_n805_), .A3(new_n866_), .A4(new_n438_), .ZN(new_n867_));
  NAND2_X1  g506(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g507(.A(new_n863_), .B1(new_n868_), .B2(G8), .ZN(new_n869_));
  INV_X1    g508(.A(new_n458_), .ZN(new_n870_));
  AOI21_X1  g509(.A(new_n457_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n871_));
  OAI21_X1  g510(.A(G8), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g511(.A1(new_n872_), .A2(KEYINPUT52), .ZN(new_n873_));
  NAND3_X1  g512(.A1(G286), .A2(new_n860_), .A3(G8), .ZN(new_n874_));
  NAND2_X1  g513(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI211_X1 g514(.A(new_n855_), .B(new_n875_), .C1(new_n865_), .C2(new_n867_), .ZN(new_n876_));
  OAI211_X1 g515(.A(new_n854_), .B(new_n859_), .C1(new_n869_), .C2(new_n876_), .ZN(new_n877_));
  INV_X1    g516(.A(G1971), .ZN(new_n878_));
  NAND2_X1  g517(.A1(new_n816_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g518(.A1(new_n819_), .A2(new_n644_), .A3(new_n809_), .ZN(new_n880_));
  NAND2_X1  g519(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g520(.A1(new_n881_), .A2(G8), .A3(G166), .ZN(new_n882_));
  NAND4_X1  g521(.A1(new_n879_), .A2(new_n880_), .A3(G8), .A4(G303), .ZN(new_n883_));
  NAND2_X1  g522(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g523(.A(KEYINPUT55), .ZN(new_n885_));
  NOR2_X1   g524(.A1(new_n816_), .A2(G2078), .ZN(new_n886_));
  OAI21_X1  g525(.A(new_n637_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n887_));
  INV_X1    g526(.A(KEYINPUT54), .ZN(new_n888_));
  NAND2_X1  g527(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g528(.A(KEYINPUT54), .B(new_n637_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n890_));
  AOI211_X1 g529(.A(new_n635_), .B(new_n886_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g530(.A1(new_n889_), .A2(new_n890_), .ZN(new_n892_));
  NAND2_X1  g531(.A1(new_n841_), .A2(new_n618_), .ZN(new_n893_));
  AOI21_X1  g532(.A(G301), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g533(.A(new_n885_), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g534(.A(new_n890_), .ZN(new_n896_));
  AOI21_X1  g535(.A(KEYINPUT54), .B1(new_n816_), .B2(new_n637_), .ZN(new_n897_));
  OAI21_X1  g536(.A(new_n893_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g537(.A1(new_n898_), .A2(new_n635_), .ZN(new_n899_));
  NAND3_X1  g538(.A1(new_n892_), .A2(G301), .A3(new_n893_), .ZN(new_n900_));
  NAND3_X1  g539(.A1(new_n899_), .A2(new_n900_), .A3(KEYINPUT55), .ZN(new_n901_));
  AOI211_X1 g540(.A(new_n877_), .B(new_n884_), .C1(new_n895_), .C2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g541(.A1(new_n846_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g542(.A1(new_n856_), .A2(new_n672_), .A3(new_n670_), .ZN(new_n904_));
  NAND4_X1  g543(.A1(new_n898_), .A2(new_n854_), .A3(new_n635_), .A4(new_n859_), .ZN(new_n905_));
  NOR2_X1   g544(.A1(new_n905_), .A2(new_n884_), .ZN(new_n906_));
  INV_X1    g545(.A(KEYINPUT61), .ZN(new_n907_));
  NAND3_X1  g546(.A1(new_n868_), .A2(G8), .A3(new_n863_), .ZN(new_n908_));
  AOI211_X1 g547(.A(new_n855_), .B(new_n863_), .C1(new_n865_), .C2(new_n867_), .ZN(new_n909_));
  OAI211_X1 g548(.A(new_n907_), .B(new_n908_), .C1(new_n909_), .C2(new_n863_), .ZN(new_n910_));
  OAI21_X1  g549(.A(KEYINPUT61), .B1(new_n869_), .B2(new_n876_), .ZN(new_n911_));
  NAND2_X1  g550(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g551(.A1(new_n906_), .A2(new_n912_), .ZN(new_n913_));
  AND2_X1   g552(.A1(new_n854_), .A2(new_n859_), .ZN(new_n914_));
  NAND4_X1  g553(.A1(new_n914_), .A2(new_n909_), .A3(new_n882_), .A4(new_n883_), .ZN(new_n915_));
  AND2_X1   g554(.A1(new_n882_), .A2(KEYINPUT62), .ZN(new_n916_));
  NOR2_X1   g555(.A1(new_n882_), .A2(KEYINPUT62), .ZN(new_n917_));
  OAI21_X1  g556(.A(new_n914_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  AND4_X1   g557(.A1(new_n904_), .A2(new_n913_), .A3(new_n915_), .A4(new_n918_), .ZN(new_n919_));
  NOR2_X1   g558(.A1(new_n841_), .A2(G288), .ZN(new_n920_));
  NAND4_X1  g559(.A1(new_n859_), .A2(G8), .A3(new_n850_), .A4(new_n920_), .ZN(new_n921_));
  NAND3_X1  g560(.A1(new_n903_), .A2(new_n919_), .A3(new_n921_), .ZN(new_n922_));
  NOR2_X1   g561(.A1(new_n819_), .A2(new_n807_), .ZN(new_n923_));
  NAND3_X1  g562(.A1(new_n923_), .A2(new_n655_), .A3(new_n653_), .ZN(new_n924_));
  NAND3_X1  g563(.A1(new_n923_), .A2(G1996), .A3(new_n748_), .ZN(new_n925_));
  AND2_X1   g564(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g565(.A1(new_n604_), .A2(G2067), .ZN(new_n927_));
  AOI21_X1  g566(.A(new_n810_), .B1(new_n597_), .B2(new_n603_), .ZN(new_n928_));
  OAI21_X1  g567(.A(new_n923_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  AND2_X1   g568(.A1(new_n926_), .A2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g569(.A1(new_n923_), .A2(new_n667_), .ZN(new_n931_));
  NOR3_X1   g570(.A1(new_n819_), .A2(new_n665_), .A3(new_n807_), .ZN(new_n932_));
  XOR2_X1   g571(.A(new_n931_), .B(new_n932_), .Z(new_n933_));
  NAND2_X1  g572(.A1(new_n930_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g573(.A1(new_n923_), .A2(G290), .ZN(new_n935_));
  XNOR2_X1  g574(.A(new_n935_), .B(KEYINPUT48), .ZN(new_n936_));
  XOR2_X1   g575(.A(KEYINPUT47), .B(G1986), .Z(new_n937_));
  NAND2_X1  g576(.A1(new_n923_), .A2(new_n937_), .ZN(new_n938_));
  AND2_X1   g577(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g578(.A1(new_n936_), .A2(new_n938_), .ZN(new_n940_));
  NOR3_X1   g579(.A1(new_n934_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g580(.A1(new_n922_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g581(.A1(new_n923_), .A2(new_n927_), .ZN(new_n943_));
  XNOR2_X1  g582(.A(new_n943_), .B(KEYINPUT50), .ZN(new_n944_));
  NOR2_X1   g583(.A1(new_n931_), .A2(new_n932_), .ZN(new_n945_));
  AOI21_X1  g584(.A(KEYINPUT49), .B1(new_n930_), .B2(new_n945_), .ZN(new_n946_));
  AOI22_X1  g585(.A1(new_n940_), .A2(new_n933_), .B1(KEYINPUT49), .B2(new_n945_), .ZN(new_n947_));
  INV_X1    g586(.A(new_n926_), .ZN(new_n948_));
  OAI21_X1  g587(.A(new_n924_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  AOI211_X1 g588(.A(new_n944_), .B(new_n946_), .C1(new_n949_), .C2(new_n929_), .ZN(new_n950_));
  NAND2_X1  g589(.A1(new_n942_), .A2(new_n950_), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g590(.A1(new_n737_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n953_));
  AOI21_X1  g591(.A(new_n769_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n954_));
  OAI21_X1  g592(.A(new_n799_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g593(.A(G227), .ZN(new_n956_));
  NAND3_X1  g594(.A1(new_n955_), .A2(KEYINPUT63), .A3(new_n956_), .ZN(new_n957_));
  INV_X1    g595(.A(KEYINPUT63), .ZN(new_n958_));
  OAI21_X1  g596(.A(new_n958_), .B1(G395), .B2(G227), .ZN(new_n959_));
  NAND2_X1  g597(.A1(new_n957_), .A2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g598(.A1(G401), .A2(G229), .ZN(new_n961_));
  AND4_X1   g599(.A1(G319), .A2(new_n960_), .A3(new_n801_), .A4(new_n961_), .ZN(G308));
  NAND4_X1  g600(.A1(new_n960_), .A2(G319), .A3(new_n801_), .A4(new_n961_), .ZN(G225));
endmodule


