//Secret key is'0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_c5315" written by ABC on Wed Oct 26 12:56:56 2022

module locked_c5315 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G4, G11, G14, G17,
    G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52,
    G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86,
    G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149,
    G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185,
    G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225,
    G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265,
    G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308,
    G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358,
    G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435,
    G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552,
    G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358,
    G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088,
    G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G4,
    G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43,
    G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81,
    G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145,
    G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179,
    G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217,
    G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257,
    G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302,
    G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348,
    G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411,
    G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545,
    G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174,
    G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087,
    G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_n384_, new_n386_, new_n396_, new_n404_, new_n405_, new_n407_,
    new_n408_, new_n412_, new_n413_, new_n414_, new_n415_, new_n417_,
    new_n418_, new_n420_, new_n421_, new_n423_, new_n424_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1007_, new_n1008_,
    new_n1010_, new_n1011_, new_n1013_, new_n1014_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1087_,
    new_n1088_, new_n1090_, new_n1091_, new_n1092_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1106_, new_n1107_, new_n1109_, new_n1110_,
    new_n1111_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1134_, new_n1135_, new_n1137_, new_n1138_, new_n1139_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1146_, new_n1147_, new_n1148_,
    new_n1150_, new_n1151_, new_n1153_, new_n1154_, new_n1155_, new_n1157_,
    new_n1158_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1208_, new_n1209_, new_n1210_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1572_, new_n1573_, new_n1574_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_;
  BUF_X1    g0000(.A(G141), .Z(G144));
  BUF_X1    g0001(.A(G293), .Z(G298));
  BUF_X1    g0002(.A(G3173), .Z(G973));
  INV_X1    g0003(.A(G545), .ZN(G594));
  INV_X1    g0004(.A(G348), .ZN(G599));
  INV_X1    g0005(.A(G366), .ZN(G600));
  INV_X1    g0006(.A(G552), .ZN(G849));
  INV_X1    g0007(.A(G562), .ZN(G850));
  NOR2_X1   g0008(.A1(G849), .A2(G850), .ZN(G601));
  INV_X1    g0009(.A(G549), .ZN(G602));
  INV_X1    g0010(.A(G545), .ZN(G603));
  INV_X1    g0011(.A(G545), .ZN(G604));
  XNOR2_X1  g0012(.A(KEYINPUT0), .B(G338), .ZN(G611));
  INV_X1    g0013(.A(G358), .ZN(G612));
  AND2_X1   g0014(.A1(G141), .A2(G145), .ZN(G810));
  INV_X1    g0015(.A(G245), .ZN(G848));
  INV_X1    g0016(.A(G559), .ZN(G851));
  AND2_X1   g0017(.A1(G1), .A2(G373), .ZN(G634));
  INV_X1    g0018(.A(G136), .ZN(new_n384_));
  NOR2_X1   g0019(.A1(new_n384_), .A2(G3173), .ZN(G815));
  INV_X1    g0020(.A(G2824), .ZN(new_n386_));
  NAND2_X1  g0021(.A1(new_n386_), .A2(G27), .ZN(G845));
  NAND2_X1  g0022(.A1(G386), .A2(G556), .ZN(G847));
  BUF_X1    g0023(.A(G137), .Z(G926));
  BUF_X1    g0024(.A(G141), .Z(G923));
  BUF_X1    g0025(.A(G1), .Z(G921));
  XNOR2_X1  g0026(.A(KEYINPUT1), .B(G549), .ZN(G892));
  BUF_X1    g0027(.A(G299), .Z(G887));
  INV_X1    g0028(.A(G549), .ZN(G606));
  NAND2_X1  g0029(.A1(G27), .A2(G31), .ZN(G809));
  INV_X1    g0030(.A(G809), .ZN(new_n396_));
  NAND2_X1  g0031(.A1(new_n396_), .A2(G140), .ZN(G656));
  BUF_X1    g0032(.A(G1), .Z(G993));
  BUF_X1    g0033(.A(G1), .Z(G978));
  BUF_X1    g0034(.A(G1), .Z(G949));
  BUF_X1    g0035(.A(G1), .Z(G939));
  BUF_X1    g0036(.A(G299), .Z(G889));
  INV_X1    g0037(.A(G299), .ZN(G593));
  INV_X1    g0038(.A(G87), .ZN(new_n404_));
  NAND2_X1  g0039(.A1(new_n404_), .A2(G2358), .ZN(new_n405_));
  OAI211_X1 g0040(.A(new_n396_), .B(new_n405_), .C1(G86), .C2(G2358), .ZN(G636));
  INV_X1    g0041(.A(G34), .ZN(new_n407_));
  NAND2_X1  g0042(.A1(new_n407_), .A2(G2358), .ZN(new_n408_));
  OAI211_X1 g0043(.A(new_n396_), .B(new_n408_), .C1(G88), .C2(G2358), .ZN(G704));
  OAI211_X1 g0044(.A(new_n396_), .B(new_n408_), .C1(G88), .C2(G2358), .ZN(G717));
  NAND2_X1  g0045(.A1(new_n396_), .A2(G83), .ZN(G820));
  INV_X1    g0046(.A(G141), .ZN(new_n412_));
  XOR2_X1   g0047(.A(KEYINPUT2), .B(G2358), .Z(new_n413_));
  NAND2_X1  g0048(.A1(new_n413_), .A2(G24), .ZN(new_n414_));
  AOI21_X1  g0049(.A(G809), .B1(G25), .B2(G2358), .ZN(new_n415_));
  AOI21_X1  g0050(.A(new_n412_), .B1(new_n414_), .B2(new_n415_), .ZN(G639));
  NAND2_X1  g0051(.A1(new_n413_), .A2(G26), .ZN(new_n417_));
  AOI21_X1  g0052(.A(G809), .B1(G81), .B2(G2358), .ZN(new_n418_));
  AOI21_X1  g0053(.A(new_n412_), .B1(new_n417_), .B2(new_n418_), .ZN(G673));
  NAND2_X1  g0054(.A1(new_n413_), .A2(G79), .ZN(new_n420_));
  AOI21_X1  g0055(.A(G809), .B1(G23), .B2(G2358), .ZN(new_n421_));
  AOI21_X1  g0056(.A(new_n412_), .B1(new_n420_), .B2(new_n421_), .ZN(G707));
  NAND2_X1  g0057(.A1(new_n413_), .A2(G82), .ZN(new_n423_));
  AOI21_X1  g0058(.A(G809), .B1(G80), .B2(G2358), .ZN(new_n424_));
  AOI21_X1  g0059(.A(new_n412_), .B1(new_n423_), .B2(new_n424_), .ZN(G715));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G341), .ZN(new_n426_));
  INV_X1    g0061(.A(G3550), .ZN(new_n427_));
  NAND2_X1  g0062(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g0063(.A(G341), .ZN(new_n429_));
  OAI211_X1 g0064(.A(new_n428_), .B(G523), .C1(new_n429_), .C2(G3552), .ZN(new_n430_));
  INV_X1    g0065(.A(new_n426_), .ZN(new_n431_));
  INV_X1    g0066(.A(G3546), .ZN(new_n432_));
  INV_X1    g0067(.A(G3548), .ZN(new_n433_));
  AOI22_X1  g0068(.A1(new_n431_), .A2(new_n432_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g0069(.A(new_n430_), .B1(new_n434_), .B2(G523), .ZN(new_n435_));
  INV_X1    g0070(.A(new_n435_), .ZN(new_n436_));
  OAI21_X1  g0071(.A(G534), .B1(G351), .B2(G3550), .ZN(new_n437_));
  INV_X1    g0072(.A(G3552), .ZN(new_n438_));
  AOI21_X1  g0073(.A(new_n437_), .B1(G351), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g0074(.A1(G351), .A2(G3546), .ZN(new_n440_));
  INV_X1    g0075(.A(G351), .ZN(new_n441_));
  AOI21_X1  g0076(.A(G534), .B1(new_n441_), .B2(G3548), .ZN(new_n442_));
  AOI21_X1  g0077(.A(new_n439_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g0078(.A(G503), .B1(G324), .B2(G3550), .ZN(new_n444_));
  AOI21_X1  g0079(.A(new_n444_), .B1(G324), .B2(new_n438_), .ZN(new_n445_));
  NAND2_X1  g0080(.A1(G324), .A2(G3546), .ZN(new_n446_));
  INV_X1    g0081(.A(G324), .ZN(new_n447_));
  AOI21_X1  g0082(.A(G503), .B1(new_n447_), .B2(G3548), .ZN(new_n448_));
  AOI21_X1  g0083(.A(new_n445_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g0084(.A1(G514), .A2(G3546), .ZN(new_n450_));
  AOI21_X1  g0085(.A(new_n450_), .B1(G514), .B2(G3552), .ZN(new_n451_));
  NAND4_X1  g0086(.A1(new_n436_), .A2(new_n443_), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  AND2_X1   g0087(.A1(new_n452_), .A2(KEYINPUT4), .ZN(new_n453_));
  NOR2_X1   g0088(.A1(new_n452_), .A2(KEYINPUT4), .ZN(new_n454_));
  NOR2_X1   g0089(.A1(G251), .A2(G302), .ZN(new_n455_));
  INV_X1    g0090(.A(G248), .ZN(new_n456_));
  AOI21_X1  g0091(.A(new_n455_), .B1(new_n456_), .B2(G302), .ZN(new_n457_));
  NOR2_X1   g0092(.A1(G251), .A2(G361), .ZN(new_n458_));
  AOI21_X1  g0093(.A(new_n458_), .B1(new_n456_), .B2(G361), .ZN(new_n459_));
  INV_X1    g0094(.A(G242), .ZN(new_n460_));
  NAND2_X1  g0095(.A1(new_n460_), .A2(G293), .ZN(new_n461_));
  OAI21_X1  g0096(.A(new_n461_), .B1(G254), .B2(G293), .ZN(new_n462_));
  NAND3_X1  g0097(.A1(new_n457_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g0098(.A1(new_n460_), .A2(G316), .ZN(new_n464_));
  INV_X1    g0099(.A(G490), .ZN(new_n465_));
  OAI211_X1 g0100(.A(new_n464_), .B(new_n465_), .C1(G254), .C2(G316), .ZN(new_n466_));
  NAND2_X1  g0101(.A1(G248), .A2(G316), .ZN(new_n467_));
  INV_X1    g0102(.A(G251), .ZN(new_n468_));
  OAI211_X1 g0103(.A(new_n467_), .B(G490), .C1(new_n468_), .C2(G316), .ZN(new_n469_));
  NAND2_X1  g0104(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g0105(.A1(new_n460_), .A2(G308), .ZN(new_n471_));
  INV_X1    g0106(.A(G479), .ZN(new_n472_));
  OAI211_X1 g0107(.A(new_n471_), .B(new_n472_), .C1(G254), .C2(G308), .ZN(new_n473_));
  NAND2_X1  g0108(.A1(G248), .A2(G308), .ZN(new_n474_));
  OAI211_X1 g0109(.A(new_n474_), .B(G479), .C1(new_n468_), .C2(G308), .ZN(new_n475_));
  NAND2_X1  g0110(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  OR3_X1    g0111(.A1(new_n463_), .A2(new_n470_), .A3(new_n476_), .ZN(new_n477_));
  NOR3_X1   g0112(.A1(new_n453_), .A2(new_n454_), .A3(new_n477_), .ZN(G598));
  NAND2_X1  g0113(.A1(G218), .A2(G468), .ZN(new_n479_));
  NOR2_X1   g0114(.A1(new_n479_), .A2(G3552), .ZN(new_n480_));
  XNOR2_X1  g0115(.A(new_n480_), .B(KEYINPUT5), .ZN(new_n481_));
  INV_X1    g0116(.A(G218), .ZN(new_n482_));
  AOI21_X1  g0117(.A(G468), .B1(new_n482_), .B2(new_n433_), .ZN(new_n483_));
  OAI21_X1  g0118(.A(new_n483_), .B1(new_n482_), .B2(G3546), .ZN(new_n484_));
  NAND2_X1  g0119(.A1(new_n482_), .A2(G468), .ZN(new_n485_));
  OAI211_X1 g0120(.A(new_n481_), .B(new_n484_), .C1(G3550), .C2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g0121(.A(new_n486_), .B(KEYINPUT6), .Z(new_n487_));
  OAI21_X1  g0122(.A(G389), .B1(G257), .B2(G3550), .ZN(new_n488_));
  AOI21_X1  g0123(.A(new_n488_), .B1(G257), .B2(new_n438_), .ZN(new_n489_));
  NAND2_X1  g0124(.A1(G257), .A2(G3546), .ZN(new_n490_));
  INV_X1    g0125(.A(G257), .ZN(new_n491_));
  AOI21_X1  g0126(.A(G389), .B1(new_n491_), .B2(G3548), .ZN(new_n492_));
  AOI21_X1  g0127(.A(new_n489_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g0128(.A1(new_n438_), .A2(G210), .A3(G457), .ZN(new_n494_));
  INV_X1    g0129(.A(G210), .ZN(new_n495_));
  NAND3_X1  g0130(.A1(new_n495_), .A2(new_n427_), .A3(G457), .ZN(new_n496_));
  INV_X1    g0131(.A(G457), .ZN(new_n497_));
  OAI21_X1  g0132(.A(new_n497_), .B1(G210), .B2(G3548), .ZN(new_n498_));
  NOR2_X1   g0133(.A1(new_n495_), .A2(G3546), .ZN(new_n499_));
  OAI211_X1 g0134(.A(new_n494_), .B(new_n496_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g0135(.A1(new_n493_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g0136(.A(G281), .ZN(new_n502_));
  AOI21_X1  g0137(.A(G374), .B1(new_n502_), .B2(G3548), .ZN(new_n503_));
  OAI21_X1  g0138(.A(new_n503_), .B1(new_n502_), .B2(new_n432_), .ZN(new_n504_));
  NOR2_X1   g0139(.A1(new_n502_), .A2(G3552), .ZN(new_n505_));
  OAI21_X1  g0140(.A(G374), .B1(G281), .B2(G3550), .ZN(new_n506_));
  OAI21_X1  g0141(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g0142(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g0143(.A1(G234), .A2(G435), .ZN(new_n509_));
  NOR2_X1   g0144(.A1(new_n509_), .A2(G3552), .ZN(new_n510_));
  XOR2_X1   g0145(.A(new_n510_), .B(KEYINPUT7), .Z(new_n511_));
  INV_X1    g0146(.A(G234), .ZN(new_n512_));
  AOI21_X1  g0147(.A(G435), .B1(new_n512_), .B2(new_n433_), .ZN(new_n513_));
  OAI21_X1  g0148(.A(new_n513_), .B1(new_n512_), .B2(G3546), .ZN(new_n514_));
  NAND2_X1  g0149(.A1(new_n512_), .A2(G435), .ZN(new_n515_));
  OAI211_X1 g0150(.A(new_n511_), .B(new_n514_), .C1(G3550), .C2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g0151(.A(G411), .B1(G273), .B2(G3550), .ZN(new_n517_));
  AOI21_X1  g0152(.A(new_n517_), .B1(G273), .B2(new_n438_), .ZN(new_n518_));
  NAND2_X1  g0153(.A1(G273), .A2(G3546), .ZN(new_n519_));
  INV_X1    g0154(.A(G273), .ZN(new_n520_));
  AOI21_X1  g0155(.A(G411), .B1(new_n520_), .B2(G3548), .ZN(new_n521_));
  AOI21_X1  g0156(.A(new_n518_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g0157(.A(new_n522_), .ZN(new_n523_));
  INV_X1    g0158(.A(G400), .ZN(new_n524_));
  OAI21_X1  g0159(.A(new_n524_), .B1(new_n433_), .B2(G265), .ZN(new_n525_));
  INV_X1    g0160(.A(G265), .ZN(new_n526_));
  NOR2_X1   g0161(.A1(new_n526_), .A2(new_n432_), .ZN(new_n527_));
  NOR2_X1   g0162(.A1(new_n526_), .A2(G3552), .ZN(new_n528_));
  OAI21_X1  g0163(.A(G400), .B1(G265), .B2(G3550), .ZN(new_n529_));
  OAI22_X1  g0164(.A1(new_n525_), .A2(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g0165(.A(G422), .ZN(new_n531_));
  OAI21_X1  g0166(.A(new_n531_), .B1(G226), .B2(G3548), .ZN(new_n532_));
  AOI21_X1  g0167(.A(new_n532_), .B1(G226), .B2(new_n432_), .ZN(new_n533_));
  INV_X1    g0168(.A(G226), .ZN(new_n534_));
  NAND3_X1  g0169(.A1(new_n534_), .A2(new_n427_), .A3(G422), .ZN(new_n535_));
  NAND2_X1  g0170(.A1(G226), .A2(G422), .ZN(new_n536_));
  OAI21_X1  g0171(.A(new_n535_), .B1(G3552), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g0172(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g0173(.A(G206), .ZN(new_n539_));
  INV_X1    g0174(.A(G254), .ZN(new_n540_));
  AOI21_X1  g0175(.A(G446), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g0176(.A(new_n541_), .B1(new_n539_), .B2(G242), .ZN(new_n542_));
  NAND2_X1  g0177(.A1(G206), .A2(G248), .ZN(new_n543_));
  OAI211_X1 g0178(.A(new_n543_), .B(G446), .C1(G206), .C2(new_n468_), .ZN(new_n544_));
  NAND2_X1  g0179(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NOR4_X1   g0180(.A1(new_n523_), .A2(new_n530_), .A3(new_n538_), .A4(new_n545_), .ZN(new_n546_));
  AND4_X1   g0181(.A1(new_n487_), .A2(new_n508_), .A3(new_n516_), .A4(new_n546_), .ZN(G610));
  INV_X1    g0182(.A(G264), .ZN(new_n548_));
  NAND2_X1  g0183(.A1(new_n548_), .A2(G335), .ZN(new_n549_));
  OAI21_X1  g0184(.A(new_n549_), .B1(G257), .B2(G335), .ZN(new_n550_));
  INV_X1    g0185(.A(G389), .ZN(new_n551_));
  NAND2_X1  g0186(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g0187(.A(new_n549_), .B(G389), .C1(G257), .C2(G335), .ZN(new_n553_));
  NAND2_X1  g0188(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g0189(.A(G335), .ZN(new_n555_));
  NOR2_X1   g0190(.A1(new_n555_), .A2(G272), .ZN(new_n556_));
  NOR2_X1   g0191(.A1(G265), .A2(G335), .ZN(new_n557_));
  OAI21_X1  g0192(.A(new_n524_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g0193(.A1(new_n526_), .A2(new_n555_), .ZN(new_n559_));
  INV_X1    g0194(.A(G272), .ZN(new_n560_));
  NAND2_X1  g0195(.A1(new_n560_), .A2(G335), .ZN(new_n561_));
  NAND3_X1  g0196(.A1(new_n559_), .A2(new_n561_), .A3(G400), .ZN(new_n562_));
  NAND2_X1  g0197(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g0198(.A1(new_n554_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g0199(.A1(new_n502_), .A2(new_n555_), .ZN(new_n565_));
  INV_X1    g0200(.A(G288), .ZN(new_n566_));
  NAND2_X1  g0201(.A1(new_n566_), .A2(G335), .ZN(new_n567_));
  NAND2_X1  g0202(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g0203(.A(G374), .ZN(new_n569_));
  NAND2_X1  g0204(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g0205(.A1(new_n565_), .A2(new_n567_), .A3(G374), .ZN(new_n571_));
  NAND2_X1  g0206(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g0207(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g0208(.A1(new_n555_), .A2(G280), .ZN(new_n574_));
  NOR2_X1   g0209(.A1(G273), .A2(G335), .ZN(new_n575_));
  NOR3_X1   g0210(.A1(new_n574_), .A2(G411), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g0211(.A(G411), .ZN(new_n577_));
  NAND2_X1  g0212(.A1(new_n520_), .A2(new_n555_), .ZN(new_n578_));
  INV_X1    g0213(.A(G280), .ZN(new_n579_));
  NAND2_X1  g0214(.A1(new_n579_), .A2(G335), .ZN(new_n580_));
  AOI21_X1  g0215(.A(new_n577_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g0216(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g0217(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g0218(.A1(new_n564_), .A2(new_n573_), .A3(new_n583_), .ZN(new_n584_));
  MUX2_X1   g0219(.A(G234), .B(G241), .S(G335), .Z(new_n585_));
  NOR2_X1   g0220(.A1(new_n585_), .A2(G435), .ZN(new_n586_));
  INV_X1    g0221(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g0222(.A1(new_n585_), .A2(G435), .ZN(new_n588_));
  NAND2_X1  g0223(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g0224(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g0225(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g0226(.A(G225), .ZN(new_n592_));
  NAND2_X1  g0227(.A1(new_n592_), .A2(G335), .ZN(new_n593_));
  OAI21_X1  g0228(.A(new_n593_), .B1(G218), .B2(G335), .ZN(new_n594_));
  INV_X1    g0229(.A(G468), .ZN(new_n595_));
  NAND2_X1  g0230(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g0231(.A(new_n593_), .B(G468), .C1(G218), .C2(G335), .ZN(new_n597_));
  AND2_X1   g0232(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g0233(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g0234(.A1(G226), .A2(G335), .ZN(new_n600_));
  INV_X1    g0235(.A(G233), .ZN(new_n601_));
  AOI21_X1  g0236(.A(new_n600_), .B1(new_n601_), .B2(G335), .ZN(new_n602_));
  NAND2_X1  g0237(.A1(new_n602_), .A2(G422), .ZN(new_n603_));
  NAND2_X1  g0238(.A1(new_n601_), .A2(G335), .ZN(new_n604_));
  OAI21_X1  g0239(.A(new_n604_), .B1(G226), .B2(G335), .ZN(new_n605_));
  NAND2_X1  g0240(.A1(new_n605_), .A2(new_n531_), .ZN(new_n606_));
  NAND2_X1  g0241(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g0242(.A1(new_n599_), .A2(new_n607_), .ZN(new_n608_));
  MUX2_X1   g0243(.A(G206), .B(G209), .S(G335), .Z(new_n609_));
  NOR2_X1   g0244(.A1(new_n609_), .A2(G446), .ZN(new_n610_));
  INV_X1    g0245(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g0246(.A1(new_n609_), .A2(G446), .ZN(new_n612_));
  NAND2_X1  g0247(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g0248(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g0249(.A1(G210), .A2(G335), .ZN(new_n615_));
  INV_X1    g0250(.A(G217), .ZN(new_n616_));
  AOI21_X1  g0251(.A(new_n615_), .B1(new_n616_), .B2(G335), .ZN(new_n617_));
  NAND2_X1  g0252(.A1(new_n617_), .A2(G457), .ZN(new_n618_));
  OR2_X1    g0253(.A1(new_n617_), .A2(G457), .ZN(new_n619_));
  NAND4_X1  g0254(.A1(new_n608_), .A2(new_n614_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n620_));
  NOR2_X1   g0255(.A1(new_n591_), .A2(new_n620_), .ZN(G588));
  INV_X1    g0256(.A(G293), .ZN(new_n622_));
  AOI21_X1  g0257(.A(G332), .B1(new_n622_), .B2(KEYINPUT8), .ZN(new_n623_));
  OAI21_X1  g0258(.A(new_n623_), .B1(KEYINPUT8), .B2(new_n622_), .ZN(new_n624_));
  NAND2_X1  g0259(.A1(G593), .A2(G332), .ZN(new_n625_));
  NAND2_X1  g0260(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g0261(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g0262(.A1(G302), .A2(G332), .ZN(new_n628_));
  INV_X1    g0263(.A(G307), .ZN(new_n629_));
  AOI21_X1  g0264(.A(new_n628_), .B1(new_n629_), .B2(G332), .ZN(new_n630_));
  NOR2_X1   g0265(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g0266(.A1(G324), .A2(G332), .ZN(new_n632_));
  INV_X1    g0267(.A(G331), .ZN(new_n633_));
  AOI21_X1  g0268(.A(new_n632_), .B1(new_n633_), .B2(G332), .ZN(new_n634_));
  AND2_X1   g0269(.A1(new_n634_), .A2(G503), .ZN(new_n635_));
  NOR2_X1   g0270(.A1(new_n634_), .A2(G503), .ZN(new_n636_));
  NOR2_X1   g0271(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g0272(.A(new_n637_), .ZN(new_n638_));
  INV_X1    g0273(.A(G332), .ZN(new_n639_));
  NOR2_X1   g0274(.A1(new_n639_), .A2(G358), .ZN(new_n640_));
  INV_X1    g0275(.A(G534), .ZN(new_n641_));
  NOR2_X1   g0276(.A1(G332), .A2(G351), .ZN(new_n642_));
  NOR3_X1   g0277(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g0278(.A1(new_n639_), .A2(new_n441_), .ZN(new_n644_));
  NAND2_X1  g0279(.A1(G612), .A2(G332), .ZN(new_n645_));
  AOI21_X1  g0280(.A(G534), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g0281(.A(KEYINPUT10), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g0282(.A(new_n641_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n648_));
  INV_X1    g0283(.A(KEYINPUT10), .ZN(new_n649_));
  NAND3_X1  g0284(.A1(new_n644_), .A2(new_n645_), .A3(G534), .ZN(new_n650_));
  NAND3_X1  g0285(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g0286(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g0287(.A(G338), .ZN(new_n653_));
  NAND2_X1  g0288(.A1(new_n653_), .A2(KEYINPUT0), .ZN(new_n654_));
  INV_X1    g0289(.A(KEYINPUT0), .ZN(new_n655_));
  NAND2_X1  g0290(.A1(new_n655_), .A2(G338), .ZN(new_n656_));
  NAND3_X1  g0291(.A1(new_n654_), .A2(new_n656_), .A3(G332), .ZN(new_n657_));
  NAND3_X1  g0292(.A1(new_n657_), .A2(KEYINPUT9), .A3(G514), .ZN(new_n658_));
  NAND2_X1  g0293(.A1(KEYINPUT9), .A2(G514), .ZN(new_n659_));
  OR2_X1    g0294(.A1(KEYINPUT9), .A2(G514), .ZN(new_n660_));
  NAND4_X1  g0295(.A1(G611), .A2(G332), .A3(new_n659_), .A4(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0296(.A1(new_n639_), .A2(new_n429_), .ZN(new_n662_));
  NAND2_X1  g0297(.A1(G599), .A2(G332), .ZN(new_n663_));
  NAND3_X1  g0298(.A1(new_n662_), .A2(new_n663_), .A3(G523), .ZN(new_n664_));
  NAND2_X1  g0299(.A1(new_n662_), .A2(new_n663_), .ZN(new_n665_));
  INV_X1    g0300(.A(G523), .ZN(new_n666_));
  NAND2_X1  g0301(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g0302(.A1(new_n658_), .A2(new_n661_), .A3(new_n664_), .A4(new_n667_), .ZN(new_n668_));
  NOR3_X1   g0303(.A1(new_n638_), .A2(new_n652_), .A3(new_n668_), .ZN(new_n669_));
  NOR2_X1   g0304(.A1(G316), .A2(G332), .ZN(new_n670_));
  INV_X1    g0305(.A(G323), .ZN(new_n671_));
  AOI21_X1  g0306(.A(new_n670_), .B1(new_n671_), .B2(G332), .ZN(new_n672_));
  NAND2_X1  g0307(.A1(new_n672_), .A2(G490), .ZN(new_n673_));
  INV_X1    g0308(.A(new_n673_), .ZN(new_n674_));
  NOR2_X1   g0309(.A1(new_n672_), .A2(G490), .ZN(new_n675_));
  NOR2_X1   g0310(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g0311(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g0312(.A1(G308), .A2(G332), .ZN(new_n678_));
  INV_X1    g0313(.A(G315), .ZN(new_n679_));
  AOI21_X1  g0314(.A(new_n678_), .B1(new_n679_), .B2(G332), .ZN(new_n680_));
  NOR2_X1   g0315(.A1(new_n680_), .A2(G479), .ZN(new_n681_));
  INV_X1    g0316(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g0317(.A1(new_n680_), .A2(G479), .ZN(new_n683_));
  NAND2_X1  g0318(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g0319(.A1(new_n677_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g0320(.A1(G600), .A2(G332), .ZN(new_n686_));
  OAI21_X1  g0321(.A(new_n686_), .B1(G332), .B2(G361), .ZN(new_n687_));
  AND4_X1   g0322(.A1(new_n631_), .A2(new_n669_), .A3(new_n685_), .A4(new_n687_), .ZN(G615));
  NOR2_X1   g0323(.A1(G332), .A2(G361), .ZN(new_n689_));
  AOI21_X1  g0324(.A(new_n689_), .B1(G332), .B2(G600), .ZN(new_n690_));
  INV_X1    g0325(.A(KEYINPUT11), .ZN(new_n691_));
  NAND2_X1  g0326(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g0327(.A1(new_n687_), .A2(KEYINPUT11), .ZN(new_n693_));
  NAND2_X1  g0328(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND4_X1   g0329(.A1(new_n631_), .A2(new_n669_), .A3(new_n685_), .A4(new_n694_), .ZN(G626));
  XOR2_X1   g0330(.A(G588), .B(KEYINPUT12), .Z(G632));
  XNOR2_X1  g0331(.A(G361), .B(G369), .ZN(new_n697_));
  XNOR2_X1  g0332(.A(new_n697_), .B(new_n447_), .ZN(new_n698_));
  XNOR2_X1  g0333(.A(G308), .B(G316), .ZN(new_n699_));
  XNOR2_X1  g0334(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g0335(.A(G341), .B(G351), .ZN(new_n701_));
  XNOR2_X1  g0336(.A(G293), .B(G302), .ZN(new_n702_));
  XNOR2_X1  g0337(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g0338(.A(new_n700_), .B(new_n703_), .ZN(G1002));
  XNOR2_X1  g0339(.A(G281), .B(G289), .ZN(new_n705_));
  XNOR2_X1  g0340(.A(new_n705_), .B(new_n512_), .ZN(new_n706_));
  AND2_X1   g0341(.A1(new_n706_), .A2(G257), .ZN(new_n707_));
  NOR2_X1   g0342(.A1(new_n706_), .A2(G257), .ZN(new_n708_));
  NOR3_X1   g0343(.A1(new_n707_), .A2(new_n708_), .A3(KEYINPUT13), .ZN(new_n709_));
  XOR2_X1   g0344(.A(G265), .B(G273), .Z(new_n710_));
  XNOR2_X1  g0345(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g0346(.A(G218), .B(G226), .ZN(new_n712_));
  XNOR2_X1  g0347(.A(G206), .B(G210), .ZN(new_n713_));
  XNOR2_X1  g0348(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g0349(.A(new_n711_), .B(new_n714_), .ZN(G1004));
  XNOR2_X1  g0350(.A(new_n597_), .B(KEYINPUT14), .ZN(new_n716_));
  NAND4_X1  g0351(.A1(new_n596_), .A2(G422), .A3(new_n597_), .A4(new_n602_), .ZN(new_n717_));
  AND2_X1   g0352(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g0353(.A1(new_n619_), .A2(new_n618_), .ZN(new_n719_));
  NOR2_X1   g0354(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g0355(.A(new_n618_), .ZN(new_n721_));
  NOR2_X1   g0356(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g0357(.A(new_n554_), .ZN(new_n723_));
  INV_X1    g0358(.A(new_n562_), .ZN(new_n724_));
  NAND2_X1  g0359(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g0360(.A1(new_n725_), .A2(new_n553_), .ZN(new_n726_));
  OAI21_X1  g0361(.A(new_n588_), .B1(new_n726_), .B2(new_n586_), .ZN(new_n727_));
  OAI211_X1 g0362(.A(new_n562_), .B(new_n558_), .C1(new_n576_), .C2(new_n581_), .ZN(new_n728_));
  INV_X1    g0363(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g0364(.A(new_n571_), .ZN(new_n730_));
  NAND2_X1  g0365(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR3_X1   g0366(.A1(new_n574_), .A2(new_n577_), .A3(new_n575_), .ZN(new_n732_));
  NAND3_X1  g0367(.A1(new_n732_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n733_));
  AOI211_X1 g0368(.A(new_n589_), .B(new_n554_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g0369(.A1(new_n727_), .A2(new_n734_), .ZN(new_n735_));
  OAI221_X1 g0370(.A(new_n612_), .B1(new_n722_), .B2(new_n610_), .C1(new_n735_), .C2(new_n620_), .ZN(G591));
  INV_X1    g0371(.A(new_n694_), .ZN(new_n737_));
  NAND2_X1  g0372(.A1(new_n669_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g0373(.A(new_n664_), .ZN(new_n739_));
  NAND3_X1  g0374(.A1(new_n658_), .A2(new_n661_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g0375(.A1(new_n657_), .A2(G514), .ZN(new_n741_));
  NAND2_X1  g0376(.A1(new_n658_), .A2(new_n661_), .ZN(new_n742_));
  NAND3_X1  g0377(.A1(new_n667_), .A2(new_n643_), .A3(new_n664_), .ZN(new_n743_));
  OAI211_X1 g0378(.A(new_n740_), .B(new_n741_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n744_));
  INV_X1    g0379(.A(new_n636_), .ZN(new_n745_));
  AOI21_X1  g0380(.A(new_n635_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g0381(.A1(new_n738_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g0382(.A1(new_n747_), .A2(new_n685_), .ZN(new_n748_));
  NAND2_X1  g0383(.A1(new_n673_), .A2(new_n683_), .ZN(new_n749_));
  NAND2_X1  g0384(.A1(new_n749_), .A2(new_n682_), .ZN(new_n750_));
  NAND3_X1  g0385(.A1(new_n748_), .A2(new_n631_), .A3(new_n750_), .ZN(G618));
  OAI221_X1 g0386(.A(new_n612_), .B1(new_n722_), .B2(new_n610_), .C1(new_n735_), .C2(new_n620_), .ZN(G621));
  NAND3_X1  g0387(.A1(new_n748_), .A2(new_n631_), .A3(new_n750_), .ZN(G629));
  INV_X1    g0388(.A(G4091), .ZN(new_n754_));
  INV_X1    g0389(.A(G4092), .ZN(new_n755_));
  OAI21_X1  g0390(.A(new_n754_), .B1(new_n755_), .B2(G131), .ZN(new_n756_));
  AOI21_X1  g0391(.A(new_n756_), .B1(new_n459_), .B2(new_n755_), .ZN(new_n757_));
  XNOR2_X1  g0392(.A(new_n687_), .B(G54), .ZN(new_n758_));
  INV_X1    g0393(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g0394(.A1(new_n754_), .A2(G4092), .ZN(new_n760_));
  AOI21_X1  g0395(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G822));
  NAND3_X1  g0396(.A1(new_n754_), .A2(G129), .A3(G4092), .ZN(new_n762_));
  XOR2_X1   g0397(.A(new_n762_), .B(KEYINPUT15), .Z(new_n763_));
  NOR2_X1   g0398(.A1(G4091), .A2(G4092), .ZN(new_n764_));
  INV_X1    g0399(.A(new_n764_), .ZN(new_n765_));
  INV_X1    g0400(.A(new_n760_), .ZN(new_n766_));
  AND3_X1   g0401(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n767_));
  AOI21_X1  g0402(.A(new_n649_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n768_));
  NOR2_X1   g0403(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g0404(.A1(new_n690_), .A2(G54), .ZN(new_n770_));
  INV_X1    g0405(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g0406(.A(new_n766_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g0407(.A(new_n772_), .ZN(new_n773_));
  NOR2_X1   g0408(.A1(new_n769_), .A2(new_n771_), .ZN(new_n774_));
  OAI221_X1 g0409(.A(new_n763_), .B1(new_n443_), .B2(new_n765_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g0410(.A(new_n775_), .ZN(G838));
  XNOR2_X1  g0411(.A(new_n572_), .B(G4), .ZN(new_n777_));
  NAND2_X1  g0412(.A1(new_n777_), .A2(new_n760_), .ZN(new_n778_));
  OR2_X1    g0413(.A1(new_n755_), .A2(G117), .ZN(new_n779_));
  OAI211_X1 g0414(.A(new_n754_), .B(new_n779_), .C1(new_n507_), .C2(G4092), .ZN(new_n780_));
  NAND2_X1  g0415(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g0416(.A(new_n781_), .ZN(G861));
  INV_X1    g0417(.A(new_n675_), .ZN(new_n783_));
  INV_X1    g0418(.A(new_n747_), .ZN(new_n784_));
  NAND3_X1  g0419(.A1(new_n669_), .A2(G54), .A3(new_n687_), .ZN(new_n785_));
  AND2_X1   g0420(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g0421(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g0422(.A(new_n783_), .B1(new_n787_), .B2(new_n674_), .ZN(new_n788_));
  AOI21_X1  g0423(.A(new_n681_), .B1(new_n788_), .B2(new_n683_), .ZN(new_n789_));
  XNOR2_X1  g0424(.A(new_n626_), .B(new_n630_), .ZN(new_n790_));
  NOR2_X1   g0425(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g0426(.A(new_n791_), .B1(new_n627_), .B2(new_n789_), .ZN(G623));
  INV_X1    g0427(.A(G822), .ZN(new_n793_));
  NOR2_X1   g0428(.A1(G4087), .A2(G4088), .ZN(new_n794_));
  NAND2_X1  g0429(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g0430(.A(G4088), .ZN(new_n796_));
  NOR2_X1   g0431(.A1(new_n796_), .A2(G61), .ZN(new_n797_));
  OAI21_X1  g0432(.A(G4087), .B1(G11), .B2(G4088), .ZN(new_n798_));
  NOR2_X1   g0433(.A1(new_n796_), .A2(G4087), .ZN(new_n799_));
  INV_X1    g0434(.A(new_n799_), .ZN(new_n800_));
  OAI221_X1 g0435(.A(new_n795_), .B1(new_n797_), .B2(new_n798_), .C1(G861), .C2(new_n800_), .ZN(G722));
  NOR2_X1   g0436(.A1(new_n652_), .A2(new_n668_), .ZN(new_n802_));
  NAND3_X1  g0437(.A1(new_n802_), .A2(G54), .A3(new_n694_), .ZN(new_n803_));
  OR2_X1    g0438(.A1(new_n742_), .A2(new_n743_), .ZN(new_n804_));
  NAND2_X1  g0439(.A1(new_n667_), .A2(new_n664_), .ZN(new_n805_));
  NOR2_X1   g0440(.A1(new_n742_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g0441(.A1(new_n806_), .A2(new_n769_), .A3(new_n690_), .ZN(new_n807_));
  NAND4_X1  g0442(.A1(new_n803_), .A2(new_n741_), .A3(new_n804_), .A4(new_n807_), .ZN(new_n808_));
  OR2_X1    g0443(.A1(new_n808_), .A2(KEYINPUT16), .ZN(new_n809_));
  NAND2_X1  g0444(.A1(new_n808_), .A2(KEYINPUT16), .ZN(new_n810_));
  NAND3_X1  g0445(.A1(new_n809_), .A2(new_n740_), .A3(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g0446(.A(new_n811_), .B(new_n638_), .ZN(new_n812_));
  AND2_X1   g0447(.A1(new_n812_), .A2(new_n760_), .ZN(new_n813_));
  OAI21_X1  g0448(.A(new_n754_), .B1(new_n755_), .B2(G52), .ZN(new_n814_));
  AOI21_X1  g0449(.A(new_n814_), .B1(new_n449_), .B2(new_n755_), .ZN(new_n815_));
  NOR2_X1   g0450(.A1(new_n813_), .A2(new_n815_), .ZN(G832));
  NAND3_X1  g0451(.A1(new_n769_), .A2(new_n667_), .A3(new_n771_), .ZN(new_n817_));
  AOI21_X1  g0452(.A(G523), .B1(new_n662_), .B2(new_n663_), .ZN(new_n818_));
  OAI21_X1  g0453(.A(new_n664_), .B1(new_n818_), .B2(new_n650_), .ZN(new_n819_));
  INV_X1    g0454(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g0455(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g0456(.A(new_n821_), .B(new_n742_), .ZN(new_n822_));
  NAND2_X1  g0457(.A1(new_n822_), .A2(new_n760_), .ZN(new_n823_));
  NAND2_X1  g0458(.A1(new_n451_), .A2(new_n755_), .ZN(new_n824_));
  OAI211_X1 g0459(.A(new_n824_), .B(new_n754_), .C1(G130), .C2(new_n755_), .ZN(new_n825_));
  NAND2_X1  g0460(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g0461(.A(new_n826_), .ZN(G834));
  NAND3_X1  g0462(.A1(new_n769_), .A2(G54), .A3(new_n694_), .ZN(new_n828_));
  OAI211_X1 g0463(.A(new_n828_), .B(new_n650_), .C1(new_n646_), .C2(new_n687_), .ZN(new_n829_));
  XNOR2_X1  g0464(.A(new_n829_), .B(new_n805_), .ZN(new_n830_));
  AND2_X1   g0465(.A1(new_n830_), .A2(new_n760_), .ZN(new_n831_));
  NOR2_X1   g0466(.A1(new_n436_), .A2(G4092), .ZN(new_n832_));
  NOR2_X1   g0467(.A1(new_n832_), .A2(KEYINPUT17), .ZN(new_n833_));
  AOI21_X1  g0468(.A(new_n833_), .B1(G119), .B2(G4092), .ZN(new_n834_));
  NAND2_X1  g0469(.A1(new_n832_), .A2(KEYINPUT17), .ZN(new_n835_));
  AOI21_X1  g0470(.A(G4091), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g0471(.A1(new_n831_), .A2(new_n836_), .ZN(G836));
  NOR2_X1   g0472(.A1(G4089), .A2(G4090), .ZN(new_n838_));
  NAND2_X1  g0473(.A1(new_n793_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g0474(.A(G4089), .ZN(new_n840_));
  NOR2_X1   g0475(.A1(new_n840_), .A2(G61), .ZN(new_n841_));
  OAI21_X1  g0476(.A(G4090), .B1(G11), .B2(G4089), .ZN(new_n842_));
  NOR2_X1   g0477(.A1(new_n840_), .A2(G4090), .ZN(new_n843_));
  INV_X1    g0478(.A(new_n843_), .ZN(new_n844_));
  OAI221_X1 g0479(.A(new_n839_), .B1(new_n841_), .B2(new_n842_), .C1(G861), .C2(new_n844_), .ZN(G859));
  INV_X1    g0480(.A(G4), .ZN(new_n846_));
  NOR2_X1   g0481(.A1(new_n572_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g0482(.A(new_n732_), .B1(new_n847_), .B2(new_n583_), .ZN(new_n848_));
  INV_X1    g0483(.A(new_n564_), .ZN(new_n849_));
  OAI22_X1  g0484(.A1(new_n848_), .A2(new_n849_), .B1(new_n731_), .B2(new_n554_), .ZN(new_n850_));
  OR2_X1    g0485(.A1(new_n850_), .A2(KEYINPUT18), .ZN(new_n851_));
  NAND2_X1  g0486(.A1(new_n850_), .A2(KEYINPUT18), .ZN(new_n852_));
  NAND3_X1  g0487(.A1(new_n851_), .A2(new_n726_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g0488(.A(new_n853_), .B(new_n589_), .ZN(new_n854_));
  NAND2_X1  g0489(.A1(new_n854_), .A2(new_n760_), .ZN(new_n855_));
  NAND2_X1  g0490(.A1(new_n516_), .A2(new_n755_), .ZN(new_n856_));
  OAI211_X1 g0491(.A(new_n856_), .B(new_n754_), .C1(G122), .C2(new_n755_), .ZN(new_n857_));
  NAND2_X1  g0492(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g0493(.A(new_n858_), .ZN(G871));
  AOI21_X1  g0494(.A(new_n724_), .B1(new_n558_), .B2(new_n732_), .ZN(new_n860_));
  NAND2_X1  g0495(.A1(new_n860_), .A2(new_n728_), .ZN(new_n861_));
  INV_X1    g0496(.A(new_n860_), .ZN(new_n862_));
  AOI21_X1  g0497(.A(G374), .B1(new_n565_), .B2(new_n567_), .ZN(new_n863_));
  OAI21_X1  g0498(.A(new_n571_), .B1(new_n863_), .B2(new_n846_), .ZN(new_n864_));
  OAI21_X1  g0499(.A(new_n861_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g0500(.A(new_n865_), .B(new_n723_), .ZN(new_n866_));
  AND2_X1   g0501(.A1(new_n866_), .A2(new_n760_), .ZN(new_n867_));
  OAI21_X1  g0502(.A(new_n754_), .B1(new_n755_), .B2(G128), .ZN(new_n868_));
  AOI21_X1  g0503(.A(new_n868_), .B1(new_n493_), .B2(new_n755_), .ZN(new_n869_));
  NOR2_X1   g0504(.A1(new_n867_), .A2(new_n869_), .ZN(G873));
  INV_X1    g0505(.A(new_n581_), .ZN(new_n871_));
  NAND3_X1  g0506(.A1(new_n578_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n872_));
  NAND3_X1  g0507(.A1(new_n871_), .A2(KEYINPUT19), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g0508(.A(KEYINPUT19), .ZN(new_n874_));
  AOI21_X1  g0509(.A(new_n571_), .B1(new_n576_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g0510(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g0511(.A1(new_n848_), .A2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g0512(.A(new_n877_), .B(new_n563_), .ZN(new_n878_));
  NAND2_X1  g0513(.A1(new_n878_), .A2(new_n760_), .ZN(new_n879_));
  OR2_X1    g0514(.A1(new_n755_), .A2(G127), .ZN(new_n880_));
  OAI211_X1 g0515(.A(new_n754_), .B(new_n880_), .C1(new_n530_), .C2(G4092), .ZN(new_n881_));
  NAND2_X1  g0516(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g0517(.A(new_n882_), .ZN(G875));
  XOR2_X1   g0518(.A(new_n864_), .B(new_n582_), .Z(new_n884_));
  NOR2_X1   g0519(.A1(new_n884_), .A2(new_n766_), .ZN(new_n885_));
  OAI21_X1  g0520(.A(new_n754_), .B1(new_n755_), .B2(G126), .ZN(new_n886_));
  AOI21_X1  g0521(.A(new_n886_), .B1(new_n522_), .B2(new_n755_), .ZN(new_n887_));
  NOR2_X1   g0522(.A1(new_n885_), .A2(new_n887_), .ZN(G877));
  MUX2_X1   g0523(.A(G369), .B(G372), .S(G332), .Z(new_n889_));
  XNOR2_X1  g0524(.A(new_n889_), .B(new_n687_), .ZN(new_n890_));
  XNOR2_X1  g0525(.A(new_n890_), .B(new_n665_), .ZN(new_n891_));
  NOR2_X1   g0526(.A1(new_n640_), .A2(new_n642_), .ZN(new_n892_));
  XNOR2_X1  g0527(.A(new_n891_), .B(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g0528(.A(new_n893_), .B(new_n790_), .ZN(new_n894_));
  NAND2_X1  g0529(.A1(new_n634_), .A2(new_n657_), .ZN(new_n895_));
  OAI21_X1  g0530(.A(new_n895_), .B1(G331), .B2(new_n657_), .ZN(new_n896_));
  XNOR2_X1  g0531(.A(new_n894_), .B(new_n896_), .ZN(new_n897_));
  INV_X1    g0532(.A(new_n680_), .ZN(new_n898_));
  XNOR2_X1  g0533(.A(new_n897_), .B(new_n898_), .ZN(new_n899_));
  XOR2_X1   g0534(.A(new_n672_), .B(KEYINPUT20), .Z(new_n900_));
  XNOR2_X1  g0535(.A(new_n899_), .B(new_n900_), .ZN(G998));
  XNOR2_X1  g0536(.A(new_n585_), .B(new_n594_), .ZN(new_n902_));
  XNOR2_X1  g0537(.A(new_n902_), .B(new_n605_), .ZN(new_n903_));
  MUX2_X1   g0538(.A(G289), .B(G292), .S(G335), .Z(new_n904_));
  XNOR2_X1  g0539(.A(new_n903_), .B(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g0540(.A(new_n550_), .B(new_n568_), .ZN(new_n906_));
  NOR2_X1   g0541(.A1(new_n574_), .A2(new_n575_), .ZN(new_n907_));
  XNOR2_X1  g0542(.A(new_n906_), .B(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g0543(.A(new_n905_), .B(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g0544(.A(new_n609_), .B(new_n617_), .ZN(new_n910_));
  NAND2_X1  g0545(.A1(new_n559_), .A2(new_n561_), .ZN(new_n911_));
  XNOR2_X1  g0546(.A(new_n910_), .B(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g0547(.A(new_n909_), .B(new_n912_), .ZN(G1000));
  NAND2_X1  g0548(.A1(new_n590_), .A2(G4), .ZN(new_n914_));
  XOR2_X1   g0549(.A(new_n914_), .B(KEYINPUT21), .Z(new_n915_));
  NAND2_X1  g0550(.A1(new_n915_), .A2(new_n735_), .ZN(new_n916_));
  AND2_X1   g0551(.A1(new_n916_), .A2(KEYINPUT22), .ZN(new_n917_));
  NOR2_X1   g0552(.A1(new_n916_), .A2(KEYINPUT22), .ZN(new_n918_));
  NOR2_X1   g0553(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g0554(.A(new_n598_), .B(new_n606_), .ZN(new_n920_));
  XNOR2_X1  g0555(.A(new_n920_), .B(KEYINPUT24), .ZN(new_n921_));
  NOR2_X1   g0556(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g0557(.A1(new_n599_), .A2(new_n603_), .ZN(new_n923_));
  NAND3_X1  g0558(.A1(new_n919_), .A2(new_n717_), .A3(new_n923_), .ZN(new_n924_));
  AOI21_X1  g0559(.A(new_n922_), .B1(KEYINPUT23), .B2(new_n924_), .ZN(new_n925_));
  OAI21_X1  g0560(.A(new_n925_), .B1(KEYINPUT23), .B2(new_n924_), .ZN(new_n926_));
  XNOR2_X1  g0561(.A(new_n722_), .B(new_n614_), .ZN(new_n927_));
  NAND2_X1  g0562(.A1(new_n919_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g0563(.A(new_n606_), .ZN(new_n929_));
  OAI21_X1  g0564(.A(new_n716_), .B1(new_n599_), .B2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g0565(.A(new_n721_), .B1(new_n930_), .B2(new_n619_), .ZN(new_n931_));
  XNOR2_X1  g0566(.A(new_n931_), .B(KEYINPUT25), .ZN(new_n932_));
  XNOR2_X1  g0567(.A(new_n932_), .B(new_n613_), .ZN(new_n933_));
  NAND2_X1  g0568(.A1(new_n933_), .A2(new_n916_), .ZN(new_n934_));
  NAND2_X1  g0569(.A1(new_n928_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g0570(.A(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g0571(.A(new_n916_), .B(new_n607_), .ZN(new_n937_));
  INV_X1    g0572(.A(new_n884_), .ZN(new_n938_));
  OR3_X1    g0573(.A1(new_n866_), .A2(new_n777_), .A3(new_n938_), .ZN(new_n939_));
  NOR4_X1   g0574(.A1(new_n937_), .A2(new_n854_), .A3(new_n878_), .A4(new_n939_), .ZN(new_n940_));
  NAND4_X1  g0575(.A1(new_n917_), .A2(new_n618_), .A3(new_n619_), .A4(new_n608_), .ZN(new_n941_));
  NAND2_X1  g0576(.A1(new_n916_), .A2(new_n608_), .ZN(new_n942_));
  NAND3_X1  g0577(.A1(new_n942_), .A2(new_n719_), .A3(new_n718_), .ZN(new_n943_));
  NOR2_X1   g0578(.A1(new_n918_), .A2(new_n720_), .ZN(new_n944_));
  NAND3_X1  g0579(.A1(new_n941_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n945_));
  INV_X1    g0580(.A(new_n945_), .ZN(new_n946_));
  OAI211_X1 g0581(.A(new_n936_), .B(new_n940_), .C1(KEYINPUT26), .C2(new_n946_), .ZN(new_n947_));
  AOI211_X1 g0582(.A(new_n926_), .B(new_n947_), .C1(KEYINPUT26), .C2(new_n946_), .ZN(G575));
  INV_X1    g0583(.A(new_n750_), .ZN(new_n949_));
  AOI21_X1  g0584(.A(new_n949_), .B1(new_n787_), .B2(new_n685_), .ZN(new_n950_));
  XNOR2_X1  g0585(.A(new_n950_), .B(new_n630_), .ZN(new_n951_));
  INV_X1    g0586(.A(new_n951_), .ZN(new_n952_));
  XNOR2_X1  g0587(.A(new_n786_), .B(new_n676_), .ZN(new_n953_));
  NOR2_X1   g0588(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  XNOR2_X1  g0589(.A(new_n788_), .B(new_n684_), .ZN(new_n955_));
  NAND3_X1  g0590(.A1(new_n954_), .A2(G623), .A3(new_n955_), .ZN(new_n956_));
  XOR2_X1   g0591(.A(new_n956_), .B(KEYINPUT27), .Z(new_n957_));
  OR3_X1    g0592(.A1(new_n830_), .A2(new_n652_), .A3(new_n759_), .ZN(new_n958_));
  NOR4_X1   g0593(.A1(new_n957_), .A2(new_n812_), .A3(new_n822_), .A4(new_n958_), .ZN(G585));
  INV_X1    g0594(.A(G137), .ZN(new_n960_));
  INV_X1    g0595(.A(G1689), .ZN(new_n961_));
  NOR2_X1   g0596(.A1(new_n961_), .A2(G1690), .ZN(new_n962_));
  NAND2_X1  g0597(.A1(new_n781_), .A2(new_n962_), .ZN(new_n963_));
  OAI21_X1  g0598(.A(G1690), .B1(G182), .B2(G1689), .ZN(new_n964_));
  INV_X1    g0599(.A(G185), .ZN(new_n965_));
  AOI21_X1  g0600(.A(new_n964_), .B1(new_n965_), .B2(G1689), .ZN(new_n966_));
  NOR2_X1   g0601(.A1(G1689), .A2(G1690), .ZN(new_n967_));
  AOI21_X1  g0602(.A(new_n966_), .B1(new_n793_), .B2(new_n967_), .ZN(new_n968_));
  AOI21_X1  g0603(.A(new_n960_), .B1(new_n963_), .B2(new_n968_), .ZN(G661));
  OR3_X1    g0604(.A1(G822), .A2(KEYINPUT28), .A3(G1694), .ZN(new_n970_));
  INV_X1    g0605(.A(G1691), .ZN(new_n971_));
  OAI21_X1  g0606(.A(KEYINPUT28), .B1(G822), .B2(G1694), .ZN(new_n972_));
  NAND3_X1  g0607(.A1(new_n970_), .A2(new_n971_), .A3(new_n972_), .ZN(new_n973_));
  OAI21_X1  g0608(.A(G1694), .B1(G182), .B2(G1691), .ZN(new_n974_));
  AOI21_X1  g0609(.A(new_n974_), .B1(new_n965_), .B2(G1691), .ZN(new_n975_));
  NOR2_X1   g0610(.A1(new_n971_), .A2(G1694), .ZN(new_n976_));
  AOI21_X1  g0611(.A(new_n975_), .B1(new_n781_), .B2(new_n976_), .ZN(new_n977_));
  AOI21_X1  g0612(.A(new_n960_), .B1(new_n973_), .B2(new_n977_), .ZN(G693));
  NAND3_X1  g0613(.A1(G37), .A2(G4087), .A3(G4088), .ZN(new_n979_));
  XNOR2_X1  g0614(.A(new_n979_), .B(KEYINPUT29), .ZN(new_n980_));
  AND3_X1   g0615(.A1(new_n796_), .A2(G43), .A3(G4087), .ZN(new_n981_));
  AOI211_X1 g0616(.A(new_n980_), .B(new_n981_), .C1(new_n858_), .C2(new_n799_), .ZN(new_n982_));
  INV_X1    g0617(.A(new_n794_), .ZN(new_n983_));
  OAI21_X1  g0618(.A(new_n982_), .B1(G832), .B2(new_n983_), .ZN(new_n984_));
  XNOR2_X1  g0619(.A(new_n984_), .B(KEYINPUT30), .ZN(G747));
  NOR2_X1   g0620(.A1(G873), .A2(new_n800_), .ZN(new_n986_));
  XNOR2_X1  g0621(.A(new_n986_), .B(KEYINPUT31), .ZN(new_n987_));
  NOR2_X1   g0622(.A1(new_n796_), .A2(G20), .ZN(new_n988_));
  OAI21_X1  g0623(.A(G4087), .B1(G76), .B2(G4088), .ZN(new_n989_));
  OAI221_X1 g0624(.A(new_n987_), .B1(new_n983_), .B2(G834), .C1(new_n988_), .C2(new_n989_), .ZN(G752));
  NAND3_X1  g0625(.A1(G17), .A2(G4087), .A3(G4088), .ZN(new_n991_));
  OR2_X1    g0626(.A1(new_n991_), .A2(KEYINPUT32), .ZN(new_n992_));
  NAND2_X1  g0627(.A1(new_n991_), .A2(KEYINPUT32), .ZN(new_n993_));
  AND2_X1   g0628(.A1(G73), .A2(G4087), .ZN(new_n994_));
  AOI22_X1  g0629(.A1(new_n992_), .A2(new_n993_), .B1(new_n796_), .B2(new_n994_), .ZN(new_n995_));
  OAI221_X1 g0630(.A(new_n995_), .B1(new_n800_), .B2(G875), .C1(G836), .C2(new_n983_), .ZN(G757));
  INV_X1    g0631(.A(G70), .ZN(new_n997_));
  NAND2_X1  g0632(.A1(new_n997_), .A2(G4088), .ZN(new_n998_));
  OAI211_X1 g0633(.A(new_n998_), .B(G4087), .C1(G67), .C2(G4088), .ZN(new_n999_));
  OAI221_X1 g0634(.A(new_n999_), .B1(new_n800_), .B2(G877), .C1(G838), .C2(new_n983_), .ZN(G762));
  NAND2_X1  g0635(.A1(new_n858_), .A2(new_n843_), .ZN(new_n1001_));
  XNOR2_X1  g0636(.A(new_n1001_), .B(KEYINPUT33), .ZN(new_n1002_));
  NOR2_X1   g0637(.A1(new_n840_), .A2(G37), .ZN(new_n1003_));
  OAI21_X1  g0638(.A(G4090), .B1(G43), .B2(G4089), .ZN(new_n1004_));
  INV_X1    g0639(.A(new_n838_), .ZN(new_n1005_));
  OAI221_X1 g0640(.A(new_n1002_), .B1(new_n1003_), .B2(new_n1004_), .C1(G832), .C2(new_n1005_), .ZN(G787));
  OR2_X1    g0641(.A1(G76), .A2(G4089), .ZN(new_n1007_));
  OAI211_X1 g0642(.A(new_n1007_), .B(G4090), .C1(G20), .C2(new_n840_), .ZN(new_n1008_));
  OAI221_X1 g0643(.A(new_n1008_), .B1(G873), .B2(new_n844_), .C1(G834), .C2(new_n1005_), .ZN(G792));
  OR2_X1    g0644(.A1(G73), .A2(G4089), .ZN(new_n1010_));
  OAI211_X1 g0645(.A(new_n1010_), .B(G4090), .C1(G17), .C2(new_n840_), .ZN(new_n1011_));
  OAI221_X1 g0646(.A(new_n1011_), .B1(new_n844_), .B2(G875), .C1(G836), .C2(new_n1005_), .ZN(G797));
  NAND2_X1  g0647(.A1(new_n997_), .A2(G4089), .ZN(new_n1013_));
  OAI211_X1 g0648(.A(new_n1013_), .B(G4090), .C1(G67), .C2(G4089), .ZN(new_n1014_));
  OAI221_X1 g0649(.A(new_n1014_), .B1(new_n844_), .B2(G877), .C1(G838), .C2(new_n1005_), .ZN(G802));
  INV_X1    g0650(.A(G832), .ZN(new_n1016_));
  NAND2_X1  g0651(.A1(new_n1016_), .A2(new_n967_), .ZN(new_n1017_));
  OAI21_X1  g0652(.A(G1690), .B1(G200), .B2(G1689), .ZN(new_n1018_));
  INV_X1    g0653(.A(G170), .ZN(new_n1019_));
  AOI21_X1  g0654(.A(new_n1018_), .B1(new_n1019_), .B2(G1689), .ZN(new_n1020_));
  AOI21_X1  g0655(.A(new_n1020_), .B1(new_n858_), .B2(new_n962_), .ZN(new_n1021_));
  AOI21_X1  g0656(.A(new_n960_), .B1(new_n1017_), .B2(new_n1021_), .ZN(G642));
  OAI21_X1  g0657(.A(G1690), .B1(G188), .B2(G1689), .ZN(new_n1023_));
  INV_X1    g0658(.A(G158), .ZN(new_n1024_));
  AOI21_X1  g0659(.A(new_n1023_), .B1(new_n1024_), .B2(G1689), .ZN(new_n1025_));
  AOI21_X1  g0660(.A(new_n1025_), .B1(new_n775_), .B2(new_n967_), .ZN(new_n1026_));
  INV_X1    g0661(.A(G877), .ZN(new_n1027_));
  NAND2_X1  g0662(.A1(new_n1027_), .A2(new_n962_), .ZN(new_n1028_));
  AOI21_X1  g0663(.A(new_n960_), .B1(new_n1026_), .B2(new_n1028_), .ZN(G664));
  OAI21_X1  g0664(.A(G1690), .B1(G155), .B2(G1689), .ZN(new_n1030_));
  INV_X1    g0665(.A(G152), .ZN(new_n1031_));
  AOI21_X1  g0666(.A(new_n1030_), .B1(new_n1031_), .B2(G1689), .ZN(new_n1032_));
  INV_X1    g0667(.A(G836), .ZN(new_n1033_));
  AOI21_X1  g0668(.A(new_n1032_), .B1(new_n1033_), .B2(new_n967_), .ZN(new_n1034_));
  NAND2_X1  g0669(.A1(new_n882_), .A2(new_n962_), .ZN(new_n1035_));
  AOI21_X1  g0670(.A(new_n960_), .B1(new_n1034_), .B2(new_n1035_), .ZN(G667));
  OAI21_X1  g0671(.A(G1690), .B1(G149), .B2(G1689), .ZN(new_n1037_));
  INV_X1    g0672(.A(G146), .ZN(new_n1038_));
  AOI21_X1  g0673(.A(new_n1037_), .B1(new_n1038_), .B2(G1689), .ZN(new_n1039_));
  AOI21_X1  g0674(.A(new_n1039_), .B1(new_n826_), .B2(new_n967_), .ZN(new_n1040_));
  INV_X1    g0675(.A(KEYINPUT34), .ZN(new_n1041_));
  OR2_X1    g0676(.A1(new_n1040_), .A2(new_n1041_), .ZN(new_n1042_));
  INV_X1    g0677(.A(G873), .ZN(new_n1043_));
  AOI22_X1  g0678(.A1(new_n1040_), .A2(new_n1041_), .B1(new_n1043_), .B2(new_n962_), .ZN(new_n1044_));
  AOI21_X1  g0679(.A(new_n960_), .B1(new_n1042_), .B2(new_n1044_), .ZN(G670));
  NOR2_X1   g0680(.A1(G1691), .A2(G1694), .ZN(new_n1046_));
  NAND2_X1  g0681(.A1(new_n1016_), .A2(new_n1046_), .ZN(new_n1047_));
  OAI21_X1  g0682(.A(G1694), .B1(G200), .B2(G1691), .ZN(new_n1048_));
  AOI21_X1  g0683(.A(new_n1048_), .B1(new_n1019_), .B2(G1691), .ZN(new_n1049_));
  AOI21_X1  g0684(.A(new_n1049_), .B1(new_n858_), .B2(new_n976_), .ZN(new_n1050_));
  AOI21_X1  g0685(.A(new_n960_), .B1(new_n1047_), .B2(new_n1050_), .ZN(G676));
  OAI21_X1  g0686(.A(G1694), .B1(G188), .B2(G1691), .ZN(new_n1052_));
  AOI21_X1  g0687(.A(new_n1052_), .B1(new_n1024_), .B2(G1691), .ZN(new_n1053_));
  AOI21_X1  g0688(.A(new_n1053_), .B1(new_n775_), .B2(new_n1046_), .ZN(new_n1054_));
  NAND2_X1  g0689(.A1(new_n1027_), .A2(new_n976_), .ZN(new_n1055_));
  AOI21_X1  g0690(.A(new_n960_), .B1(new_n1054_), .B2(new_n1055_), .ZN(G696));
  NAND2_X1  g0691(.A1(new_n1031_), .A2(G1691), .ZN(new_n1057_));
  OAI211_X1 g0692(.A(new_n1057_), .B(G1694), .C1(G155), .C2(G1691), .ZN(new_n1058_));
  INV_X1    g0693(.A(new_n976_), .ZN(new_n1059_));
  INV_X1    g0694(.A(new_n1046_), .ZN(new_n1060_));
  OAI221_X1 g0695(.A(new_n1058_), .B1(G875), .B2(new_n1059_), .C1(G836), .C2(new_n1060_), .ZN(new_n1061_));
  NAND2_X1  g0696(.A1(new_n1061_), .A2(G137), .ZN(new_n1062_));
  XOR2_X1   g0697(.A(new_n1062_), .B(KEYINPUT35), .Z(G699));
  NOR2_X1   g0698(.A1(G834), .A2(G1694), .ZN(new_n1064_));
  AOI21_X1  g0699(.A(G1691), .B1(new_n1064_), .B2(KEYINPUT37), .ZN(new_n1065_));
  OAI21_X1  g0700(.A(new_n1065_), .B1(KEYINPUT37), .B2(new_n1064_), .ZN(new_n1066_));
  NAND3_X1  g0701(.A1(G146), .A2(G1691), .A3(G1694), .ZN(new_n1067_));
  NOR2_X1   g0702(.A1(new_n1067_), .A2(KEYINPUT36), .ZN(new_n1068_));
  NAND2_X1  g0703(.A1(new_n1067_), .A2(KEYINPUT36), .ZN(new_n1069_));
  NAND3_X1  g0704(.A1(new_n971_), .A2(G149), .A3(G1694), .ZN(new_n1070_));
  NAND2_X1  g0705(.A1(new_n1069_), .A2(new_n1070_), .ZN(new_n1071_));
  AOI211_X1 g0706(.A(new_n1068_), .B(new_n1071_), .C1(new_n1043_), .C2(new_n976_), .ZN(new_n1072_));
  AOI21_X1  g0707(.A(new_n960_), .B1(new_n1066_), .B2(new_n1072_), .ZN(G702));
  NAND2_X1  g0708(.A1(G135), .A2(G4115), .ZN(new_n1074_));
  NOR2_X1   g0709(.A1(new_n462_), .A2(G3717), .ZN(new_n1075_));
  INV_X1    g0710(.A(G3724), .ZN(new_n1076_));
  INV_X1    g0711(.A(G123), .ZN(new_n1077_));
  INV_X1    g0712(.A(G3717), .ZN(new_n1078_));
  OAI21_X1  g0713(.A(new_n1076_), .B1(new_n1077_), .B2(new_n1078_), .ZN(new_n1079_));
  OAI21_X1  g0714(.A(new_n1074_), .B1(new_n1075_), .B2(new_n1079_), .ZN(new_n1080_));
  INV_X1    g0715(.A(G623), .ZN(new_n1081_));
  NAND2_X1  g0716(.A1(new_n1081_), .A2(G3717), .ZN(new_n1082_));
  XOR2_X1   g0717(.A(new_n626_), .B(G132), .Z(new_n1083_));
  AOI21_X1  g0718(.A(new_n1076_), .B1(new_n1083_), .B2(new_n1078_), .ZN(new_n1084_));
  AOI21_X1  g0719(.A(new_n1080_), .B1(new_n1082_), .B2(new_n1084_), .ZN(G818));
  XNOR2_X1  g0720(.A(G623), .B(new_n1083_), .ZN(G813));
  OAI21_X1  g0721(.A(new_n754_), .B1(new_n755_), .B2(G123), .ZN(new_n1087_));
  AOI21_X1  g0722(.A(new_n1087_), .B1(new_n462_), .B2(new_n755_), .ZN(new_n1088_));
  AOI21_X1  g0723(.A(new_n1088_), .B1(new_n1081_), .B2(new_n760_), .ZN(G824));
  OAI21_X1  g0724(.A(new_n754_), .B1(new_n755_), .B2(G121), .ZN(new_n1090_));
  AOI21_X1  g0725(.A(new_n1090_), .B1(new_n457_), .B2(new_n755_), .ZN(new_n1091_));
  AOI21_X1  g0726(.A(new_n1091_), .B1(new_n952_), .B2(new_n760_), .ZN(new_n1092_));
  XNOR2_X1  g0727(.A(new_n1092_), .B(KEYINPUT38), .ZN(G826));
  AOI21_X1  g0728(.A(G4092), .B1(new_n473_), .B2(new_n475_), .ZN(new_n1094_));
  NAND2_X1  g0729(.A1(G116), .A2(G4092), .ZN(new_n1095_));
  XNOR2_X1  g0730(.A(new_n1095_), .B(KEYINPUT39), .ZN(new_n1096_));
  OAI21_X1  g0731(.A(new_n754_), .B1(new_n1094_), .B2(new_n1096_), .ZN(new_n1097_));
  XNOR2_X1  g0732(.A(new_n1097_), .B(KEYINPUT40), .ZN(new_n1098_));
  OAI21_X1  g0733(.A(new_n1098_), .B1(new_n955_), .B2(new_n766_), .ZN(new_n1099_));
  INV_X1    g0734(.A(new_n1099_), .ZN(G828));
  NAND2_X1  g0735(.A1(new_n953_), .A2(new_n760_), .ZN(new_n1101_));
  OR2_X1    g0736(.A1(new_n755_), .A2(G112), .ZN(new_n1102_));
  OAI211_X1 g0737(.A(new_n754_), .B(new_n1102_), .C1(new_n470_), .C2(G4092), .ZN(new_n1103_));
  NAND2_X1  g0738(.A1(new_n1101_), .A2(new_n1103_), .ZN(new_n1104_));
  INV_X1    g0739(.A(new_n1104_), .ZN(G830));
  NAND3_X1  g0740(.A1(G601), .A2(G245), .A3(G559), .ZN(new_n1106_));
  OR3_X1    g0741(.A1(G1002), .A2(G847), .A3(new_n1106_), .ZN(new_n1107_));
  NOR4_X1   g0742(.A1(G998), .A2(G1004), .A3(G1000), .A4(new_n1107_), .ZN(G854));
  OAI21_X1  g0743(.A(new_n754_), .B1(new_n755_), .B2(G115), .ZN(new_n1109_));
  INV_X1    g0744(.A(new_n545_), .ZN(new_n1110_));
  AOI21_X1  g0745(.A(new_n1109_), .B1(new_n1110_), .B2(new_n755_), .ZN(new_n1111_));
  AOI21_X1  g0746(.A(new_n1111_), .B1(new_n935_), .B2(new_n760_), .ZN(G863));
  NAND2_X1  g0747(.A1(new_n500_), .A2(new_n755_), .ZN(new_n1113_));
  OAI211_X1 g0748(.A(new_n1113_), .B(new_n754_), .C1(G114), .C2(new_n755_), .ZN(new_n1114_));
  OAI21_X1  g0749(.A(new_n1114_), .B1(new_n945_), .B2(new_n766_), .ZN(new_n1115_));
  XNOR2_X1  g0750(.A(new_n1115_), .B(KEYINPUT41), .ZN(new_n1116_));
  INV_X1    g0751(.A(new_n1116_), .ZN(G865));
  AND2_X1   g0752(.A1(new_n926_), .A2(new_n760_), .ZN(new_n1118_));
  AND2_X1   g0753(.A1(new_n1118_), .A2(KEYINPUT42), .ZN(new_n1119_));
  NAND2_X1  g0754(.A1(new_n487_), .A2(new_n755_), .ZN(new_n1120_));
  OAI211_X1 g0755(.A(new_n1120_), .B(new_n754_), .C1(G53), .C2(new_n755_), .ZN(new_n1121_));
  OAI21_X1  g0756(.A(new_n1121_), .B1(new_n1118_), .B2(KEYINPUT42), .ZN(new_n1122_));
  NOR2_X1   g0757(.A1(new_n1119_), .A2(new_n1122_), .ZN(G867));
  AND2_X1   g0758(.A1(new_n937_), .A2(new_n760_), .ZN(new_n1124_));
  OAI21_X1  g0759(.A(new_n754_), .B1(new_n755_), .B2(G113), .ZN(new_n1125_));
  INV_X1    g0760(.A(new_n538_), .ZN(new_n1126_));
  AOI21_X1  g0761(.A(new_n1125_), .B1(new_n1126_), .B2(new_n755_), .ZN(new_n1127_));
  NOR2_X1   g0762(.A1(new_n1124_), .A2(new_n1127_), .ZN(G869));
  INV_X1    g0763(.A(G106), .ZN(new_n1129_));
  NAND2_X1  g0764(.A1(new_n1129_), .A2(G4089), .ZN(new_n1130_));
  OAI211_X1 g0765(.A(new_n1130_), .B(G4090), .C1(G109), .C2(G4089), .ZN(new_n1131_));
  XNOR2_X1  g0766(.A(G863), .B(KEYINPUT43), .ZN(new_n1132_));
  OAI221_X1 g0767(.A(new_n1131_), .B1(new_n1005_), .B2(G824), .C1(new_n1132_), .C2(new_n844_), .ZN(G712));
  NAND2_X1  g0768(.A1(new_n1129_), .A2(G4088), .ZN(new_n1134_));
  OAI211_X1 g0769(.A(new_n1134_), .B(G4087), .C1(G109), .C2(G4088), .ZN(new_n1135_));
  OAI221_X1 g0770(.A(new_n1135_), .B1(new_n983_), .B2(G824), .C1(new_n1132_), .C2(new_n800_), .ZN(G727));
  INV_X1    g0771(.A(G49), .ZN(new_n1137_));
  NAND2_X1  g0772(.A1(new_n1137_), .A2(G4088), .ZN(new_n1138_));
  OAI211_X1 g0773(.A(new_n1138_), .B(G4087), .C1(G46), .C2(G4088), .ZN(new_n1139_));
  OAI221_X1 g0774(.A(new_n1139_), .B1(G826), .B2(new_n983_), .C1(G865), .C2(new_n800_), .ZN(G732));
  OAI21_X1  g0775(.A(G4087), .B1(G100), .B2(G4088), .ZN(new_n1141_));
  INV_X1    g0776(.A(G103), .ZN(new_n1142_));
  AOI21_X1  g0777(.A(new_n1141_), .B1(new_n1142_), .B2(G4088), .ZN(new_n1143_));
  AOI21_X1  g0778(.A(new_n1143_), .B1(new_n1099_), .B2(new_n794_), .ZN(new_n1144_));
  OAI21_X1  g0779(.A(new_n1144_), .B1(G867), .B2(new_n800_), .ZN(G737));
  INV_X1    g0780(.A(G40), .ZN(new_n1146_));
  NAND2_X1  g0781(.A1(new_n1146_), .A2(G4088), .ZN(new_n1147_));
  OAI211_X1 g0782(.A(new_n1147_), .B(G4087), .C1(G91), .C2(G4088), .ZN(new_n1148_));
  OAI221_X1 g0783(.A(new_n1148_), .B1(new_n983_), .B2(G830), .C1(G869), .C2(new_n800_), .ZN(G742));
  NAND2_X1  g0784(.A1(new_n1137_), .A2(G4089), .ZN(new_n1150_));
  OAI211_X1 g0785(.A(new_n1150_), .B(G4090), .C1(G46), .C2(G4089), .ZN(new_n1151_));
  OAI221_X1 g0786(.A(new_n1151_), .B1(G826), .B2(new_n1005_), .C1(G865), .C2(new_n844_), .ZN(G772));
  OAI21_X1  g0787(.A(G4090), .B1(G100), .B2(G4089), .ZN(new_n1153_));
  AOI21_X1  g0788(.A(new_n1153_), .B1(new_n1142_), .B2(G4089), .ZN(new_n1154_));
  AOI21_X1  g0789(.A(new_n1154_), .B1(new_n1099_), .B2(new_n838_), .ZN(new_n1155_));
  OAI21_X1  g0790(.A(new_n1155_), .B1(G867), .B2(new_n844_), .ZN(G777));
  NAND2_X1  g0791(.A1(new_n1146_), .A2(G4089), .ZN(new_n1157_));
  OAI211_X1 g0792(.A(new_n1157_), .B(G4090), .C1(G91), .C2(G4089), .ZN(new_n1158_));
  OAI221_X1 g0793(.A(new_n1158_), .B1(new_n1005_), .B2(G830), .C1(G869), .C2(new_n844_), .ZN(G782));
  NAND3_X1  g0794(.A1(G173), .A2(G1689), .A3(G1690), .ZN(new_n1160_));
  OR2_X1    g0795(.A1(new_n1160_), .A2(KEYINPUT44), .ZN(new_n1161_));
  NAND2_X1  g0796(.A1(new_n1160_), .A2(KEYINPUT44), .ZN(new_n1162_));
  AOI21_X1  g0797(.A(KEYINPUT45), .B1(G203), .B2(G1690), .ZN(new_n1163_));
  NAND3_X1  g0798(.A1(KEYINPUT45), .A2(G203), .A3(G1690), .ZN(new_n1164_));
  NAND2_X1  g0799(.A1(new_n1164_), .A2(new_n961_), .ZN(new_n1165_));
  OAI211_X1 g0800(.A(new_n1161_), .B(new_n1162_), .C1(new_n1163_), .C2(new_n1165_), .ZN(new_n1166_));
  INV_X1    g0801(.A(G869), .ZN(new_n1167_));
  AOI21_X1  g0802(.A(new_n1166_), .B1(new_n1167_), .B2(new_n962_), .ZN(new_n1168_));
  NAND2_X1  g0803(.A1(new_n1104_), .A2(new_n967_), .ZN(new_n1169_));
  AOI21_X1  g0804(.A(new_n960_), .B1(new_n1168_), .B2(new_n1169_), .ZN(G645));
  INV_X1    g0805(.A(G867), .ZN(new_n1171_));
  NAND2_X1  g0806(.A1(new_n1171_), .A2(new_n962_), .ZN(new_n1172_));
  OAI21_X1  g0807(.A(G1690), .B1(G197), .B2(G1689), .ZN(new_n1173_));
  INV_X1    g0808(.A(G167), .ZN(new_n1174_));
  AOI21_X1  g0809(.A(new_n1173_), .B1(new_n1174_), .B2(G1689), .ZN(new_n1175_));
  AOI21_X1  g0810(.A(new_n1175_), .B1(new_n1099_), .B2(new_n967_), .ZN(new_n1176_));
  AOI21_X1  g0811(.A(new_n960_), .B1(new_n1172_), .B2(new_n1176_), .ZN(G648));
  INV_X1    g0812(.A(G826), .ZN(new_n1178_));
  NAND2_X1  g0813(.A1(new_n1178_), .A2(new_n967_), .ZN(new_n1179_));
  OAI21_X1  g0814(.A(G1690), .B1(G194), .B2(G1689), .ZN(new_n1180_));
  INV_X1    g0815(.A(G164), .ZN(new_n1181_));
  AOI21_X1  g0816(.A(new_n1180_), .B1(new_n1181_), .B2(G1689), .ZN(new_n1182_));
  AOI21_X1  g0817(.A(new_n1182_), .B1(new_n1116_), .B2(new_n962_), .ZN(new_n1183_));
  AOI21_X1  g0818(.A(new_n960_), .B1(new_n1179_), .B2(new_n1183_), .ZN(G651));
  INV_X1    g0819(.A(G161), .ZN(new_n1185_));
  NAND2_X1  g0820(.A1(new_n1185_), .A2(G1689), .ZN(new_n1186_));
  OAI211_X1 g0821(.A(new_n1186_), .B(G1690), .C1(G191), .C2(G1689), .ZN(new_n1187_));
  INV_X1    g0822(.A(new_n967_), .ZN(new_n1188_));
  INV_X1    g0823(.A(new_n962_), .ZN(new_n1189_));
  OAI221_X1 g0824(.A(new_n1187_), .B1(new_n1188_), .B2(G824), .C1(new_n1132_), .C2(new_n1189_), .ZN(new_n1190_));
  AND2_X1   g0825(.A1(new_n1190_), .A2(G137), .ZN(G654));
  OAI21_X1  g0826(.A(G1694), .B1(G203), .B2(G1691), .ZN(new_n1192_));
  INV_X1    g0827(.A(G173), .ZN(new_n1193_));
  AOI21_X1  g0828(.A(new_n1192_), .B1(new_n1193_), .B2(G1691), .ZN(new_n1194_));
  AOI21_X1  g0829(.A(new_n1194_), .B1(new_n1167_), .B2(new_n976_), .ZN(new_n1195_));
  NAND2_X1  g0830(.A1(new_n1104_), .A2(new_n1046_), .ZN(new_n1196_));
  AOI21_X1  g0831(.A(new_n960_), .B1(new_n1195_), .B2(new_n1196_), .ZN(G679));
  NAND2_X1  g0832(.A1(new_n1171_), .A2(new_n976_), .ZN(new_n1198_));
  OAI21_X1  g0833(.A(G1694), .B1(G197), .B2(G1691), .ZN(new_n1199_));
  AOI21_X1  g0834(.A(new_n1199_), .B1(new_n1174_), .B2(G1691), .ZN(new_n1200_));
  AOI21_X1  g0835(.A(new_n1200_), .B1(new_n1099_), .B2(new_n1046_), .ZN(new_n1201_));
  AOI21_X1  g0836(.A(new_n960_), .B1(new_n1198_), .B2(new_n1201_), .ZN(G682));
  NAND2_X1  g0837(.A1(new_n1178_), .A2(new_n1046_), .ZN(new_n1203_));
  OAI21_X1  g0838(.A(G1694), .B1(G194), .B2(G1691), .ZN(new_n1204_));
  AOI21_X1  g0839(.A(new_n1204_), .B1(new_n1181_), .B2(G1691), .ZN(new_n1205_));
  AOI21_X1  g0840(.A(new_n1205_), .B1(new_n1116_), .B2(new_n976_), .ZN(new_n1206_));
  AOI21_X1  g0841(.A(new_n960_), .B1(new_n1203_), .B2(new_n1206_), .ZN(G685));
  NAND2_X1  g0842(.A1(new_n1185_), .A2(G1691), .ZN(new_n1208_));
  OAI211_X1 g0843(.A(new_n1208_), .B(G1694), .C1(G191), .C2(G1691), .ZN(new_n1209_));
  OAI221_X1 g0844(.A(new_n1209_), .B1(new_n1060_), .B2(G824), .C1(new_n1132_), .C2(new_n1059_), .ZN(new_n1210_));
  AND2_X1   g0845(.A1(new_n1210_), .A2(G137), .ZN(G688));
  AOI21_X1  g0846(.A(new_n641_), .B1(G251), .B2(new_n441_), .ZN(new_n1212_));
  OAI21_X1  g0847(.A(new_n1212_), .B1(new_n456_), .B2(new_n441_), .ZN(new_n1213_));
  AOI21_X1  g0848(.A(G534), .B1(new_n540_), .B2(new_n441_), .ZN(new_n1214_));
  OAI21_X1  g0849(.A(new_n1214_), .B1(G242), .B2(new_n441_), .ZN(new_n1215_));
  NAND2_X1  g0850(.A1(new_n1213_), .A2(new_n1215_), .ZN(new_n1216_));
  XNOR2_X1  g0851(.A(new_n1216_), .B(new_n459_), .ZN(new_n1217_));
  MUX2_X1   g0852(.A(new_n460_), .B(G248), .S(G514), .Z(new_n1218_));
  XNOR2_X1  g0853(.A(new_n1217_), .B(new_n1218_), .ZN(new_n1219_));
  XNOR2_X1  g0854(.A(new_n457_), .B(new_n462_), .ZN(new_n1220_));
  XNOR2_X1  g0855(.A(new_n1219_), .B(new_n1220_), .ZN(new_n1221_));
  AOI21_X1  g0856(.A(G523), .B1(new_n429_), .B2(G254), .ZN(new_n1222_));
  OAI21_X1  g0857(.A(new_n1222_), .B1(new_n460_), .B2(new_n429_), .ZN(new_n1223_));
  AOI22_X1  g0858(.A1(new_n426_), .A2(G251), .B1(G248), .B2(G341), .ZN(new_n1224_));
  OAI21_X1  g0859(.A(new_n1223_), .B1(new_n1224_), .B2(new_n666_), .ZN(new_n1225_));
  NAND2_X1  g0860(.A1(G248), .A2(G324), .ZN(new_n1226_));
  INV_X1    g0861(.A(G503), .ZN(new_n1227_));
  AOI21_X1  g0862(.A(new_n1227_), .B1(G251), .B2(new_n447_), .ZN(new_n1228_));
  AOI21_X1  g0863(.A(G503), .B1(new_n540_), .B2(new_n447_), .ZN(new_n1229_));
  NAND2_X1  g0864(.A1(new_n460_), .A2(G324), .ZN(new_n1230_));
  AOI22_X1  g0865(.A1(new_n1226_), .A2(new_n1228_), .B1(new_n1229_), .B2(new_n1230_), .ZN(new_n1231_));
  XNOR2_X1  g0866(.A(new_n1225_), .B(new_n1231_), .ZN(new_n1232_));
  XNOR2_X1  g0867(.A(new_n470_), .B(new_n476_), .ZN(new_n1233_));
  XNOR2_X1  g0868(.A(new_n1232_), .B(new_n1233_), .ZN(new_n1234_));
  XNOR2_X1  g0869(.A(new_n1221_), .B(new_n1234_), .ZN(new_n1235_));
  NAND2_X1  g0870(.A1(new_n1235_), .A2(new_n764_), .ZN(new_n1236_));
  OAI21_X1  g0871(.A(G4092), .B1(G120), .B2(G4091), .ZN(new_n1237_));
  NAND3_X1  g0872(.A1(new_n669_), .A2(G2174), .A3(new_n694_), .ZN(new_n1238_));
  NAND2_X1  g0873(.A1(new_n784_), .A2(new_n1238_), .ZN(new_n1239_));
  OAI21_X1  g0874(.A(new_n749_), .B1(new_n673_), .B2(new_n681_), .ZN(new_n1240_));
  OAI21_X1  g0875(.A(new_n1240_), .B1(new_n949_), .B2(new_n630_), .ZN(new_n1241_));
  NOR4_X1   g0876(.A1(new_n673_), .A2(G479), .A3(new_n630_), .A4(new_n680_), .ZN(new_n1242_));
  INV_X1    g0877(.A(KEYINPUT54), .ZN(new_n1243_));
  OR2_X1    g0878(.A1(new_n1242_), .A2(new_n1243_), .ZN(new_n1244_));
  NAND2_X1  g0879(.A1(new_n1242_), .A2(new_n1243_), .ZN(new_n1245_));
  NAND3_X1  g0880(.A1(new_n1241_), .A2(new_n1244_), .A3(new_n1245_), .ZN(new_n1246_));
  NAND2_X1  g0881(.A1(new_n1246_), .A2(new_n677_), .ZN(new_n1247_));
  INV_X1    g0882(.A(new_n684_), .ZN(new_n1248_));
  INV_X1    g0883(.A(new_n630_), .ZN(new_n1249_));
  NAND2_X1  g0884(.A1(new_n676_), .A2(new_n1249_), .ZN(new_n1250_));
  NAND3_X1  g0885(.A1(new_n1247_), .A2(new_n1248_), .A3(new_n1250_), .ZN(new_n1251_));
  NAND2_X1  g0886(.A1(new_n1251_), .A2(KEYINPUT55), .ZN(new_n1252_));
  INV_X1    g0887(.A(KEYINPUT55), .ZN(new_n1253_));
  NAND4_X1  g0888(.A1(new_n1247_), .A2(new_n1253_), .A3(new_n1248_), .A4(new_n1250_), .ZN(new_n1254_));
  NAND2_X1  g0889(.A1(new_n1246_), .A2(new_n676_), .ZN(new_n1255_));
  NOR2_X1   g0890(.A1(new_n1242_), .A2(new_n676_), .ZN(new_n1256_));
  AOI21_X1  g0891(.A(new_n1248_), .B1(new_n1241_), .B2(new_n1256_), .ZN(new_n1257_));
  NAND2_X1  g0892(.A1(new_n1255_), .A2(new_n1257_), .ZN(new_n1258_));
  NAND3_X1  g0893(.A1(new_n1252_), .A2(new_n1254_), .A3(new_n1258_), .ZN(new_n1259_));
  XNOR2_X1  g0894(.A(new_n1259_), .B(new_n630_), .ZN(new_n1260_));
  AOI21_X1  g0895(.A(new_n1239_), .B1(new_n1260_), .B2(new_n626_), .ZN(new_n1261_));
  OAI21_X1  g0896(.A(new_n1261_), .B1(new_n626_), .B2(new_n1260_), .ZN(new_n1262_));
  NAND2_X1  g0897(.A1(new_n898_), .A2(new_n630_), .ZN(new_n1263_));
  XNOR2_X1  g0898(.A(new_n1263_), .B(new_n675_), .ZN(new_n1264_));
  OAI21_X1  g0899(.A(new_n1264_), .B1(new_n1249_), .B2(new_n684_), .ZN(new_n1265_));
  AOI21_X1  g0900(.A(KEYINPUT53), .B1(new_n1265_), .B2(new_n676_), .ZN(new_n1266_));
  XNOR2_X1  g0901(.A(new_n684_), .B(new_n626_), .ZN(new_n1267_));
  NOR2_X1   g0902(.A1(new_n1266_), .A2(new_n1267_), .ZN(new_n1268_));
  XNOR2_X1  g0903(.A(new_n676_), .B(new_n630_), .ZN(new_n1269_));
  XNOR2_X1  g0904(.A(new_n1265_), .B(new_n1269_), .ZN(new_n1270_));
  XNOR2_X1  g0905(.A(new_n1268_), .B(new_n1270_), .ZN(new_n1271_));
  NAND2_X1  g0906(.A1(new_n1271_), .A2(new_n1239_), .ZN(new_n1272_));
  NAND2_X1  g0907(.A1(new_n1262_), .A2(new_n1272_), .ZN(new_n1273_));
  INV_X1    g0908(.A(new_n1273_), .ZN(new_n1274_));
  NAND2_X1  g0909(.A1(new_n648_), .A2(new_n650_), .ZN(new_n1275_));
  OAI211_X1 g0910(.A(new_n743_), .B(new_n664_), .C1(new_n1275_), .C2(new_n818_), .ZN(new_n1276_));
  AOI22_X1  g0911(.A1(new_n1276_), .A2(new_n690_), .B1(new_n694_), .B2(new_n820_), .ZN(new_n1277_));
  NAND3_X1  g0912(.A1(new_n647_), .A2(new_n651_), .A3(new_n690_), .ZN(new_n1278_));
  INV_X1    g0913(.A(KEYINPUT47), .ZN(new_n1279_));
  AND3_X1   g0914(.A1(new_n1278_), .A2(new_n1279_), .A3(new_n650_), .ZN(new_n1280_));
  AOI21_X1  g0915(.A(new_n1279_), .B1(new_n1278_), .B2(new_n650_), .ZN(new_n1281_));
  OAI21_X1  g0916(.A(new_n1277_), .B1(new_n1280_), .B2(new_n1281_), .ZN(new_n1282_));
  NAND2_X1  g0917(.A1(new_n1278_), .A2(new_n650_), .ZN(new_n1283_));
  NAND2_X1  g0918(.A1(new_n1283_), .A2(KEYINPUT47), .ZN(new_n1284_));
  NOR2_X1   g0919(.A1(new_n1275_), .A2(new_n818_), .ZN(new_n1285_));
  OAI21_X1  g0920(.A(new_n690_), .B1(new_n1285_), .B2(new_n819_), .ZN(new_n1286_));
  NAND2_X1  g0921(.A1(new_n820_), .A2(new_n694_), .ZN(new_n1287_));
  NAND2_X1  g0922(.A1(new_n1286_), .A2(new_n1287_), .ZN(new_n1288_));
  NAND3_X1  g0923(.A1(new_n1278_), .A2(new_n1279_), .A3(new_n650_), .ZN(new_n1289_));
  NAND3_X1  g0924(.A1(new_n1284_), .A2(new_n1288_), .A3(new_n1289_), .ZN(new_n1290_));
  NAND3_X1  g0925(.A1(new_n1282_), .A2(new_n1290_), .A3(KEYINPUT48), .ZN(new_n1291_));
  NOR3_X1   g0926(.A1(new_n652_), .A2(new_n668_), .A3(new_n687_), .ZN(new_n1292_));
  OAI21_X1  g0927(.A(KEYINPUT46), .B1(new_n1292_), .B2(new_n744_), .ZN(new_n1293_));
  INV_X1    g0928(.A(new_n744_), .ZN(new_n1294_));
  INV_X1    g0929(.A(KEYINPUT46), .ZN(new_n1295_));
  NAND3_X1  g0930(.A1(new_n1294_), .A2(new_n807_), .A3(new_n1295_), .ZN(new_n1296_));
  NAND2_X1  g0931(.A1(new_n1293_), .A2(new_n1296_), .ZN(new_n1297_));
  NAND2_X1  g0932(.A1(new_n1284_), .A2(new_n1289_), .ZN(new_n1298_));
  INV_X1    g0933(.A(KEYINPUT48), .ZN(new_n1299_));
  NAND3_X1  g0934(.A1(new_n1298_), .A2(new_n1299_), .A3(new_n1277_), .ZN(new_n1300_));
  AND3_X1   g0935(.A1(new_n1291_), .A2(new_n1297_), .A3(new_n1300_), .ZN(new_n1301_));
  NAND2_X1  g0936(.A1(new_n1276_), .A2(new_n737_), .ZN(new_n1302_));
  NAND2_X1  g0937(.A1(new_n820_), .A2(new_n687_), .ZN(new_n1303_));
  AND2_X1   g0938(.A1(new_n1302_), .A2(new_n1303_), .ZN(new_n1304_));
  OAI21_X1  g0939(.A(new_n648_), .B1(new_n737_), .B2(new_n643_), .ZN(new_n1305_));
  OAI21_X1  g0940(.A(new_n1282_), .B1(new_n1304_), .B2(new_n1305_), .ZN(new_n1306_));
  OAI21_X1  g0941(.A(new_n690_), .B1(new_n1306_), .B2(new_n1297_), .ZN(new_n1307_));
  OAI21_X1  g0942(.A(KEYINPUT49), .B1(new_n1301_), .B2(new_n1307_), .ZN(new_n1308_));
  NOR3_X1   g0943(.A1(new_n1292_), .A2(KEYINPUT46), .A3(new_n744_), .ZN(new_n1309_));
  AOI21_X1  g0944(.A(new_n1295_), .B1(new_n1294_), .B2(new_n807_), .ZN(new_n1310_));
  NOR2_X1   g0945(.A1(new_n1309_), .A2(new_n1310_), .ZN(new_n1311_));
  NAND3_X1  g0946(.A1(new_n1291_), .A2(new_n1311_), .A3(new_n1300_), .ZN(new_n1312_));
  AOI21_X1  g0947(.A(new_n1305_), .B1(new_n1302_), .B2(new_n1303_), .ZN(new_n1313_));
  AOI21_X1  g0948(.A(new_n1313_), .B1(new_n1298_), .B2(new_n1277_), .ZN(new_n1314_));
  NAND2_X1  g0949(.A1(new_n1314_), .A2(new_n1297_), .ZN(new_n1315_));
  NAND3_X1  g0950(.A1(new_n1312_), .A2(new_n694_), .A3(new_n1315_), .ZN(new_n1316_));
  AOI21_X1  g0951(.A(new_n687_), .B1(new_n1314_), .B2(new_n1311_), .ZN(new_n1317_));
  NAND3_X1  g0952(.A1(new_n1291_), .A2(new_n1297_), .A3(new_n1300_), .ZN(new_n1318_));
  INV_X1    g0953(.A(KEYINPUT49), .ZN(new_n1319_));
  NAND3_X1  g0954(.A1(new_n1317_), .A2(new_n1318_), .A3(new_n1319_), .ZN(new_n1320_));
  NAND4_X1  g0955(.A1(new_n1308_), .A2(new_n652_), .A3(new_n1316_), .A4(new_n1320_), .ZN(new_n1321_));
  AND3_X1   g0956(.A1(new_n1312_), .A2(new_n694_), .A3(new_n1315_), .ZN(new_n1322_));
  AOI21_X1  g0957(.A(new_n694_), .B1(new_n1312_), .B2(new_n1315_), .ZN(new_n1323_));
  OAI21_X1  g0958(.A(new_n769_), .B1(new_n1322_), .B2(new_n1323_), .ZN(new_n1324_));
  NAND3_X1  g0959(.A1(new_n1321_), .A2(new_n1324_), .A3(new_n638_), .ZN(new_n1325_));
  INV_X1    g0960(.A(KEYINPUT50), .ZN(new_n1326_));
  NAND2_X1  g0961(.A1(new_n1325_), .A2(new_n1326_), .ZN(new_n1327_));
  NAND4_X1  g0962(.A1(new_n1308_), .A2(new_n769_), .A3(new_n1316_), .A4(new_n1320_), .ZN(new_n1328_));
  OAI21_X1  g0963(.A(new_n652_), .B1(new_n1322_), .B2(new_n1323_), .ZN(new_n1329_));
  NAND3_X1  g0964(.A1(new_n1328_), .A2(new_n1329_), .A3(new_n637_), .ZN(new_n1330_));
  NAND4_X1  g0965(.A1(new_n1321_), .A2(new_n1324_), .A3(KEYINPUT50), .A4(new_n638_), .ZN(new_n1331_));
  NAND3_X1  g0966(.A1(new_n1327_), .A2(new_n1330_), .A3(new_n1331_), .ZN(new_n1332_));
  NAND2_X1  g0967(.A1(new_n742_), .A2(new_n805_), .ZN(new_n1333_));
  AND2_X1   g0968(.A1(new_n1333_), .A2(new_n668_), .ZN(new_n1334_));
  INV_X1    g0969(.A(new_n1334_), .ZN(new_n1335_));
  NAND2_X1  g0970(.A1(new_n1332_), .A2(new_n1335_), .ZN(new_n1336_));
  AND2_X1   g0971(.A1(new_n1330_), .A2(new_n1334_), .ZN(new_n1337_));
  NAND2_X1  g0972(.A1(new_n1328_), .A2(new_n1329_), .ZN(new_n1338_));
  NAND2_X1  g0973(.A1(new_n1338_), .A2(new_n638_), .ZN(new_n1339_));
  NAND2_X1  g0974(.A1(new_n1337_), .A2(new_n1339_), .ZN(new_n1340_));
  AOI21_X1  g0975(.A(G2174), .B1(new_n1336_), .B2(new_n1340_), .ZN(new_n1341_));
  INV_X1    g0976(.A(G2174), .ZN(new_n1342_));
  XNOR2_X1  g0977(.A(new_n637_), .B(new_n694_), .ZN(new_n1343_));
  XNOR2_X1  g0978(.A(new_n1343_), .B(new_n1334_), .ZN(new_n1344_));
  INV_X1    g0979(.A(new_n1344_), .ZN(new_n1345_));
  AOI211_X1 g0980(.A(new_n643_), .B(new_n820_), .C1(new_n648_), .C2(new_n692_), .ZN(new_n1346_));
  XOR2_X1   g0981(.A(new_n1346_), .B(KEYINPUT51), .Z(new_n1347_));
  OAI21_X1  g0982(.A(new_n1298_), .B1(new_n1275_), .B2(new_n690_), .ZN(new_n1348_));
  AOI21_X1  g0983(.A(new_n819_), .B1(new_n1285_), .B2(new_n692_), .ZN(new_n1349_));
  NAND2_X1  g0984(.A1(new_n1348_), .A2(new_n1349_), .ZN(new_n1350_));
  INV_X1    g0985(.A(KEYINPUT52), .ZN(new_n1351_));
  NAND2_X1  g0986(.A1(new_n802_), .A2(new_n694_), .ZN(new_n1352_));
  NAND3_X1  g0987(.A1(new_n1352_), .A2(new_n1294_), .A3(new_n807_), .ZN(new_n1353_));
  OAI211_X1 g0988(.A(new_n1347_), .B(new_n1350_), .C1(new_n1351_), .C2(new_n1353_), .ZN(new_n1354_));
  NAND2_X1  g0989(.A1(new_n1353_), .A2(new_n1351_), .ZN(new_n1355_));
  XNOR2_X1  g0990(.A(new_n1354_), .B(new_n1355_), .ZN(new_n1356_));
  OR2_X1    g0991(.A1(new_n1356_), .A2(new_n652_), .ZN(new_n1357_));
  OAI21_X1  g0992(.A(new_n1356_), .B1(new_n691_), .B2(new_n652_), .ZN(new_n1358_));
  AOI21_X1  g0993(.A(new_n1345_), .B1(new_n1357_), .B2(new_n1358_), .ZN(new_n1359_));
  INV_X1    g0994(.A(new_n1359_), .ZN(new_n1360_));
  NAND3_X1  g0995(.A1(new_n1357_), .A2(new_n1358_), .A3(new_n1345_), .ZN(new_n1361_));
  AOI21_X1  g0996(.A(new_n1342_), .B1(new_n1360_), .B2(new_n1361_), .ZN(new_n1362_));
  OAI21_X1  g0997(.A(new_n1274_), .B1(new_n1341_), .B2(new_n1362_), .ZN(new_n1363_));
  INV_X1    g0998(.A(new_n1361_), .ZN(new_n1364_));
  OAI21_X1  g0999(.A(G2174), .B1(new_n1364_), .B2(new_n1359_), .ZN(new_n1365_));
  AOI22_X1  g1000(.A1(new_n1332_), .A2(new_n1335_), .B1(new_n1339_), .B2(new_n1337_), .ZN(new_n1366_));
  OAI211_X1 g1001(.A(new_n1365_), .B(new_n1273_), .C1(new_n1366_), .C2(G2174), .ZN(new_n1367_));
  NAND2_X1  g1002(.A1(new_n1363_), .A2(new_n1367_), .ZN(new_n1368_));
  OAI211_X1 g1003(.A(new_n1236_), .B(new_n1237_), .C1(new_n1368_), .C2(new_n766_), .ZN(G843));
  XNOR2_X1  g1004(.A(new_n598_), .B(new_n607_), .ZN(new_n1370_));
  MUX2_X1   g1005(.A(new_n597_), .B(new_n596_), .S(new_n606_), .Z(new_n1371_));
  MUX2_X1   g1006(.A(new_n607_), .B(new_n1370_), .S(new_n1371_), .Z(new_n1372_));
  XNOR2_X1  g1007(.A(new_n1372_), .B(new_n931_), .ZN(new_n1373_));
  XOR2_X1   g1008(.A(new_n613_), .B(new_n719_), .Z(new_n1374_));
  INV_X1    g1009(.A(new_n1374_), .ZN(new_n1375_));
  OR2_X1    g1010(.A1(new_n1373_), .A2(new_n1375_), .ZN(new_n1376_));
  NAND2_X1  g1011(.A1(new_n1373_), .A2(new_n1375_), .ZN(new_n1377_));
  NAND3_X1  g1012(.A1(new_n735_), .A2(G1497), .A3(new_n591_), .ZN(new_n1378_));
  INV_X1    g1013(.A(new_n1378_), .ZN(new_n1379_));
  NOR3_X1   g1014(.A1(new_n727_), .A2(new_n734_), .A3(G1497), .ZN(new_n1380_));
  NOR2_X1   g1015(.A1(new_n1379_), .A2(new_n1380_), .ZN(new_n1381_));
  NAND3_X1  g1016(.A1(new_n1376_), .A2(new_n1377_), .A3(new_n1381_), .ZN(new_n1382_));
  INV_X1    g1017(.A(new_n1382_), .ZN(new_n1383_));
  MUX2_X1   g1018(.A(new_n596_), .B(new_n597_), .S(new_n603_), .Z(new_n1384_));
  MUX2_X1   g1019(.A(new_n607_), .B(new_n1370_), .S(new_n1384_), .Z(new_n1385_));
  XNOR2_X1  g1020(.A(new_n1385_), .B(new_n722_), .ZN(new_n1386_));
  NOR2_X1   g1021(.A1(new_n599_), .A2(KEYINPUT56), .ZN(new_n1387_));
  NAND2_X1  g1022(.A1(new_n1386_), .A2(new_n1387_), .ZN(new_n1388_));
  INV_X1    g1023(.A(new_n1388_), .ZN(new_n1389_));
  INV_X1    g1024(.A(KEYINPUT56), .ZN(new_n1390_));
  NOR2_X1   g1025(.A1(new_n1386_), .A2(new_n1390_), .ZN(new_n1391_));
  OAI21_X1  g1026(.A(new_n1374_), .B1(new_n1389_), .B2(new_n1391_), .ZN(new_n1392_));
  OAI211_X1 g1027(.A(new_n1388_), .B(new_n1375_), .C1(new_n1390_), .C2(new_n1386_), .ZN(new_n1393_));
  NAND2_X1  g1028(.A1(new_n1392_), .A2(new_n1393_), .ZN(new_n1394_));
  AOI21_X1  g1029(.A(new_n1383_), .B1(new_n1394_), .B2(new_n1380_), .ZN(new_n1395_));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1396_));
  AOI21_X1  g1031(.A(new_n1396_), .B1(new_n1394_), .B2(new_n1379_), .ZN(new_n1397_));
  AOI211_X1 g1032(.A(KEYINPUT57), .B(new_n1378_), .C1(new_n1392_), .C2(new_n1393_), .ZN(new_n1398_));
  OAI21_X1  g1033(.A(new_n1395_), .B1(new_n1397_), .B2(new_n1398_), .ZN(new_n1399_));
  AOI21_X1  g1034(.A(new_n863_), .B1(new_n860_), .B2(new_n728_), .ZN(new_n1400_));
  NAND2_X1  g1035(.A1(new_n907_), .A2(G411), .ZN(new_n1401_));
  AOI21_X1  g1036(.A(G400), .B1(new_n559_), .B2(new_n561_), .ZN(new_n1402_));
  OAI211_X1 g1037(.A(new_n863_), .B(new_n562_), .C1(new_n1401_), .C2(new_n1402_), .ZN(new_n1403_));
  INV_X1    g1038(.A(new_n1403_), .ZN(new_n1404_));
  OAI21_X1  g1039(.A(KEYINPUT59), .B1(new_n1400_), .B2(new_n1404_), .ZN(new_n1405_));
  OAI211_X1 g1040(.A(new_n570_), .B(new_n571_), .C1(new_n576_), .C2(new_n581_), .ZN(new_n1406_));
  AOI21_X1  g1041(.A(new_n732_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n1407_));
  NAND3_X1  g1042(.A1(new_n1405_), .A2(new_n1406_), .A3(new_n1407_), .ZN(new_n1408_));
  NAND2_X1  g1043(.A1(new_n1407_), .A2(new_n1406_), .ZN(new_n1409_));
  OAI211_X1 g1044(.A(new_n1409_), .B(KEYINPUT59), .C1(new_n1400_), .C2(new_n1404_), .ZN(new_n1410_));
  OAI211_X1 g1045(.A(new_n733_), .B(new_n553_), .C1(new_n728_), .C2(new_n571_), .ZN(new_n1411_));
  NAND2_X1  g1046(.A1(new_n1411_), .A2(new_n552_), .ZN(new_n1412_));
  NAND2_X1  g1047(.A1(new_n1412_), .A2(new_n584_), .ZN(new_n1413_));
  INV_X1    g1048(.A(KEYINPUT58), .ZN(new_n1414_));
  OAI21_X1  g1049(.A(new_n725_), .B1(new_n1413_), .B2(new_n1414_), .ZN(new_n1415_));
  NOR3_X1   g1050(.A1(new_n1406_), .A2(new_n554_), .A3(new_n563_), .ZN(new_n1416_));
  AOI21_X1  g1051(.A(new_n1416_), .B1(new_n552_), .B2(new_n1411_), .ZN(new_n1417_));
  NOR2_X1   g1052(.A1(new_n1417_), .A2(KEYINPUT58), .ZN(new_n1418_));
  OAI211_X1 g1053(.A(new_n1408_), .B(new_n1410_), .C1(new_n1415_), .C2(new_n1418_), .ZN(new_n1419_));
  AOI22_X1  g1054(.A1(new_n1417_), .A2(KEYINPUT58), .B1(new_n723_), .B2(new_n724_), .ZN(new_n1420_));
  NOR2_X1   g1055(.A1(new_n1400_), .A2(new_n1404_), .ZN(new_n1421_));
  NAND2_X1  g1056(.A1(new_n1421_), .A2(new_n1409_), .ZN(new_n1422_));
  OAI211_X1 g1057(.A(new_n1406_), .B(new_n1407_), .C1(new_n1400_), .C2(new_n1404_), .ZN(new_n1423_));
  NAND2_X1  g1058(.A1(new_n1413_), .A2(new_n1414_), .ZN(new_n1424_));
  NAND4_X1  g1059(.A1(new_n1420_), .A2(new_n1422_), .A3(new_n1423_), .A4(new_n1424_), .ZN(new_n1425_));
  AND3_X1   g1060(.A1(new_n1419_), .A2(new_n1425_), .A3(new_n572_), .ZN(new_n1426_));
  AOI21_X1  g1061(.A(new_n572_), .B1(new_n1419_), .B2(new_n1425_), .ZN(new_n1427_));
  OAI21_X1  g1062(.A(new_n582_), .B1(new_n1426_), .B2(new_n1427_), .ZN(new_n1428_));
  INV_X1    g1063(.A(new_n589_), .ZN(new_n1429_));
  NAND2_X1  g1064(.A1(new_n1408_), .A2(new_n1410_), .ZN(new_n1430_));
  AOI21_X1  g1065(.A(new_n1430_), .B1(new_n1424_), .B2(new_n1420_), .ZN(new_n1431_));
  NAND2_X1  g1066(.A1(new_n1422_), .A2(new_n1423_), .ZN(new_n1432_));
  NOR3_X1   g1067(.A1(new_n1415_), .A2(new_n1432_), .A3(new_n1418_), .ZN(new_n1433_));
  OAI21_X1  g1068(.A(new_n573_), .B1(new_n1431_), .B2(new_n1433_), .ZN(new_n1434_));
  NAND3_X1  g1069(.A1(new_n1430_), .A2(new_n1424_), .A3(new_n1420_), .ZN(new_n1435_));
  OAI21_X1  g1070(.A(new_n1432_), .B1(new_n1415_), .B2(new_n1418_), .ZN(new_n1436_));
  NAND3_X1  g1071(.A1(new_n1435_), .A2(new_n1436_), .A3(new_n572_), .ZN(new_n1437_));
  NAND3_X1  g1072(.A1(new_n1434_), .A2(new_n583_), .A3(new_n1437_), .ZN(new_n1438_));
  NAND3_X1  g1073(.A1(new_n1428_), .A2(new_n1429_), .A3(new_n1438_), .ZN(new_n1439_));
  OAI21_X1  g1074(.A(new_n583_), .B1(new_n1426_), .B2(new_n1427_), .ZN(new_n1440_));
  NAND3_X1  g1075(.A1(new_n1434_), .A2(new_n582_), .A3(new_n1437_), .ZN(new_n1441_));
  NAND3_X1  g1076(.A1(new_n1440_), .A2(new_n589_), .A3(new_n1441_), .ZN(new_n1442_));
  NAND2_X1  g1077(.A1(new_n1439_), .A2(new_n1442_), .ZN(new_n1443_));
  INV_X1    g1078(.A(new_n563_), .ZN(new_n1444_));
  OAI21_X1  g1079(.A(new_n554_), .B1(new_n1443_), .B2(new_n1444_), .ZN(new_n1445_));
  NAND2_X1  g1080(.A1(new_n1428_), .A2(new_n1438_), .ZN(new_n1446_));
  NAND2_X1  g1081(.A1(new_n1446_), .A2(new_n589_), .ZN(new_n1447_));
  AOI21_X1  g1082(.A(new_n563_), .B1(new_n1447_), .B2(new_n1439_), .ZN(new_n1448_));
  NOR2_X1   g1083(.A1(new_n1445_), .A2(new_n1448_), .ZN(new_n1449_));
  NAND2_X1  g1084(.A1(new_n1443_), .A2(new_n1444_), .ZN(new_n1450_));
  NAND3_X1  g1085(.A1(new_n1447_), .A2(new_n563_), .A3(new_n1439_), .ZN(new_n1451_));
  AOI21_X1  g1086(.A(new_n554_), .B1(new_n1450_), .B2(new_n1451_), .ZN(new_n1452_));
  OAI21_X1  g1087(.A(G1497), .B1(new_n1449_), .B2(new_n1452_), .ZN(new_n1453_));
  NAND2_X1  g1088(.A1(new_n582_), .A2(new_n572_), .ZN(new_n1454_));
  NAND2_X1  g1089(.A1(new_n1454_), .A2(new_n1406_), .ZN(new_n1455_));
  INV_X1    g1090(.A(new_n1407_), .ZN(new_n1456_));
  AOI21_X1  g1091(.A(new_n1456_), .B1(new_n1412_), .B2(new_n725_), .ZN(new_n1457_));
  INV_X1    g1092(.A(new_n1457_), .ZN(new_n1458_));
  NAND3_X1  g1093(.A1(new_n1412_), .A2(new_n725_), .A3(new_n1456_), .ZN(new_n1459_));
  AOI21_X1  g1094(.A(new_n1455_), .B1(new_n1458_), .B2(new_n1459_), .ZN(new_n1460_));
  INV_X1    g1095(.A(new_n1459_), .ZN(new_n1461_));
  INV_X1    g1096(.A(new_n1455_), .ZN(new_n1462_));
  NOR3_X1   g1097(.A1(new_n1461_), .A2(new_n1457_), .A3(new_n1462_), .ZN(new_n1463_));
  OAI21_X1  g1098(.A(new_n558_), .B1(new_n1456_), .B2(new_n724_), .ZN(new_n1464_));
  AND2_X1   g1099(.A1(new_n1464_), .A2(new_n730_), .ZN(new_n1465_));
  NOR2_X1   g1100(.A1(new_n860_), .A2(new_n730_), .ZN(new_n1466_));
  OAI22_X1  g1101(.A1(new_n1460_), .A2(new_n1463_), .B1(new_n1465_), .B2(new_n1466_), .ZN(new_n1467_));
  OAI21_X1  g1102(.A(new_n1462_), .B1(new_n1461_), .B2(new_n1457_), .ZN(new_n1468_));
  NAND3_X1  g1103(.A1(new_n1458_), .A2(new_n1459_), .A3(new_n1455_), .ZN(new_n1469_));
  AOI21_X1  g1104(.A(new_n1466_), .B1(new_n1464_), .B2(new_n730_), .ZN(new_n1470_));
  NAND3_X1  g1105(.A1(new_n1468_), .A2(new_n1469_), .A3(new_n1470_), .ZN(new_n1471_));
  NAND3_X1  g1106(.A1(new_n1467_), .A2(new_n589_), .A3(new_n1471_), .ZN(new_n1472_));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1473_));
  AOI21_X1  g1108(.A(new_n1444_), .B1(new_n1472_), .B2(new_n1473_), .ZN(new_n1474_));
  INV_X1    g1109(.A(new_n1471_), .ZN(new_n1475_));
  AOI21_X1  g1110(.A(new_n1470_), .B1(new_n1468_), .B2(new_n1469_), .ZN(new_n1476_));
  OAI21_X1  g1111(.A(new_n1429_), .B1(new_n1475_), .B2(new_n1476_), .ZN(new_n1477_));
  NAND2_X1  g1112(.A1(new_n1477_), .A2(new_n1472_), .ZN(new_n1478_));
  NAND2_X1  g1113(.A1(new_n1474_), .A2(new_n1478_), .ZN(new_n1479_));
  OAI211_X1 g1114(.A(new_n1477_), .B(new_n1472_), .C1(new_n1473_), .C2(new_n1444_), .ZN(new_n1480_));
  NAND2_X1  g1115(.A1(new_n1479_), .A2(new_n1480_), .ZN(new_n1481_));
  NAND2_X1  g1116(.A1(new_n1481_), .A2(new_n554_), .ZN(new_n1482_));
  INV_X1    g1117(.A(G1497), .ZN(new_n1483_));
  NAND3_X1  g1118(.A1(new_n1479_), .A2(new_n723_), .A3(new_n1480_), .ZN(new_n1484_));
  NAND3_X1  g1119(.A1(new_n1482_), .A2(new_n1483_), .A3(new_n1484_), .ZN(new_n1485_));
  AOI21_X1  g1120(.A(new_n1399_), .B1(new_n1453_), .B2(new_n1485_), .ZN(new_n1486_));
  NAND2_X1  g1121(.A1(new_n1485_), .A2(new_n1399_), .ZN(new_n1487_));
  INV_X1    g1122(.A(new_n1439_), .ZN(new_n1488_));
  AOI21_X1  g1123(.A(new_n1429_), .B1(new_n1428_), .B2(new_n1438_), .ZN(new_n1489_));
  NOR3_X1   g1124(.A1(new_n1488_), .A2(new_n1444_), .A3(new_n1489_), .ZN(new_n1490_));
  AOI21_X1  g1125(.A(new_n563_), .B1(new_n1439_), .B2(new_n1442_), .ZN(new_n1491_));
  OAI21_X1  g1126(.A(new_n723_), .B1(new_n1490_), .B2(new_n1491_), .ZN(new_n1492_));
  NAND3_X1  g1127(.A1(new_n1450_), .A2(new_n1451_), .A3(new_n554_), .ZN(new_n1493_));
  NAND2_X1  g1128(.A1(new_n1492_), .A2(new_n1493_), .ZN(new_n1494_));
  AOI21_X1  g1129(.A(new_n1487_), .B1(new_n1494_), .B2(G1497), .ZN(new_n1495_));
  OAI21_X1  g1130(.A(new_n760_), .B1(new_n1486_), .B2(new_n1495_), .ZN(new_n1496_));
  OAI21_X1  g1131(.A(G4092), .B1(G118), .B2(G4091), .ZN(new_n1497_));
  AOI21_X1  g1132(.A(new_n569_), .B1(G251), .B2(new_n502_), .ZN(new_n1498_));
  OAI21_X1  g1133(.A(new_n1498_), .B1(new_n456_), .B2(new_n502_), .ZN(new_n1499_));
  AOI21_X1  g1134(.A(G374), .B1(new_n540_), .B2(new_n502_), .ZN(new_n1500_));
  OAI21_X1  g1135(.A(new_n1500_), .B1(G242), .B2(new_n502_), .ZN(new_n1501_));
  NAND2_X1  g1136(.A1(new_n1499_), .A2(new_n1501_), .ZN(new_n1502_));
  AOI21_X1  g1137(.A(new_n524_), .B1(G251), .B2(new_n526_), .ZN(new_n1503_));
  OAI21_X1  g1138(.A(new_n1503_), .B1(new_n456_), .B2(new_n526_), .ZN(new_n1504_));
  AOI21_X1  g1139(.A(G400), .B1(new_n540_), .B2(new_n526_), .ZN(new_n1505_));
  OAI21_X1  g1140(.A(new_n1505_), .B1(G242), .B2(new_n526_), .ZN(new_n1506_));
  NAND2_X1  g1141(.A1(new_n1504_), .A2(new_n1506_), .ZN(new_n1507_));
  XOR2_X1   g1142(.A(new_n1502_), .B(new_n1507_), .Z(new_n1508_));
  AOI21_X1  g1143(.A(G435), .B1(new_n512_), .B2(G254), .ZN(new_n1509_));
  OAI21_X1  g1144(.A(new_n1509_), .B1(new_n512_), .B2(new_n460_), .ZN(new_n1510_));
  OAI221_X1 g1145(.A(new_n1510_), .B1(new_n456_), .B2(new_n509_), .C1(new_n468_), .C2(new_n515_), .ZN(new_n1511_));
  XNOR2_X1  g1146(.A(new_n1508_), .B(new_n1511_), .ZN(new_n1512_));
  OAI21_X1  g1147(.A(new_n551_), .B1(new_n460_), .B2(new_n491_), .ZN(new_n1513_));
  OR2_X1    g1148(.A1(new_n1513_), .A2(KEYINPUT61), .ZN(new_n1514_));
  NAND2_X1  g1149(.A1(new_n1513_), .A2(KEYINPUT61), .ZN(new_n1515_));
  OAI211_X1 g1150(.A(new_n1514_), .B(new_n1515_), .C1(new_n540_), .C2(G257), .ZN(new_n1516_));
  NOR2_X1   g1151(.A1(new_n491_), .A2(G248), .ZN(new_n1517_));
  OAI21_X1  g1152(.A(G389), .B1(G251), .B2(G257), .ZN(new_n1518_));
  OAI21_X1  g1153(.A(new_n1516_), .B1(new_n1517_), .B2(new_n1518_), .ZN(new_n1519_));
  NAND2_X1  g1154(.A1(G248), .A2(G273), .ZN(new_n1520_));
  AOI21_X1  g1155(.A(new_n577_), .B1(G251), .B2(new_n520_), .ZN(new_n1521_));
  AOI21_X1  g1156(.A(G411), .B1(new_n540_), .B2(new_n520_), .ZN(new_n1522_));
  NAND2_X1  g1157(.A1(new_n460_), .A2(G273), .ZN(new_n1523_));
  AOI22_X1  g1158(.A1(new_n1520_), .A2(new_n1521_), .B1(new_n1522_), .B2(new_n1523_), .ZN(new_n1524_));
  XNOR2_X1  g1159(.A(new_n1519_), .B(new_n1524_), .ZN(new_n1525_));
  XNOR2_X1  g1160(.A(new_n1512_), .B(new_n1525_), .ZN(new_n1526_));
  AOI21_X1  g1161(.A(G468), .B1(new_n482_), .B2(G254), .ZN(new_n1527_));
  OAI21_X1  g1162(.A(new_n1527_), .B1(new_n482_), .B2(new_n460_), .ZN(new_n1528_));
  OAI221_X1 g1163(.A(new_n1528_), .B1(new_n456_), .B2(new_n479_), .C1(new_n468_), .C2(new_n485_), .ZN(new_n1529_));
  XNOR2_X1  g1164(.A(new_n1529_), .B(new_n545_), .ZN(new_n1530_));
  NOR2_X1   g1165(.A1(new_n536_), .A2(new_n456_), .ZN(new_n1531_));
  NOR3_X1   g1166(.A1(new_n468_), .A2(new_n531_), .A3(G226), .ZN(new_n1532_));
  NAND2_X1  g1167(.A1(G226), .A2(G242), .ZN(new_n1533_));
  AOI21_X1  g1168(.A(G422), .B1(new_n534_), .B2(G254), .ZN(new_n1534_));
  AOI211_X1 g1169(.A(new_n1531_), .B(new_n1532_), .C1(new_n1533_), .C2(new_n1534_), .ZN(new_n1535_));
  XNOR2_X1  g1170(.A(new_n1530_), .B(new_n1535_), .ZN(new_n1536_));
  XNOR2_X1  g1171(.A(new_n1526_), .B(new_n1536_), .ZN(new_n1537_));
  NOR3_X1   g1172(.A1(new_n468_), .A2(new_n497_), .A3(G210), .ZN(new_n1538_));
  NOR3_X1   g1173(.A1(new_n495_), .A2(new_n456_), .A3(new_n497_), .ZN(new_n1539_));
  NAND2_X1  g1174(.A1(G210), .A2(G242), .ZN(new_n1540_));
  AOI21_X1  g1175(.A(G457), .B1(new_n495_), .B2(G254), .ZN(new_n1541_));
  AOI211_X1 g1176(.A(new_n1538_), .B(new_n1539_), .C1(new_n1540_), .C2(new_n1541_), .ZN(new_n1542_));
  AOI21_X1  g1177(.A(new_n765_), .B1(new_n1537_), .B2(new_n1542_), .ZN(new_n1543_));
  OAI21_X1  g1178(.A(new_n1543_), .B1(new_n1542_), .B2(new_n1537_), .ZN(new_n1544_));
  XNOR2_X1  g1179(.A(new_n1544_), .B(KEYINPUT62), .ZN(new_n1545_));
  NAND3_X1  g1180(.A1(new_n1496_), .A2(new_n1497_), .A3(new_n1545_), .ZN(G882));
  OAI21_X1  g1181(.A(G4087), .B1(G14), .B2(G4088), .ZN(new_n1547_));
  INV_X1    g1182(.A(G64), .ZN(new_n1548_));
  AOI21_X1  g1183(.A(new_n1547_), .B1(new_n1548_), .B2(G4088), .ZN(new_n1549_));
  OR2_X1    g1184(.A1(new_n755_), .A2(G97), .ZN(new_n1550_));
  NAND2_X1  g1185(.A1(new_n1544_), .A2(new_n1550_), .ZN(new_n1551_));
  INV_X1    g1186(.A(new_n1399_), .ZN(new_n1552_));
  OAI21_X1  g1187(.A(new_n1444_), .B1(new_n1488_), .B2(new_n1489_), .ZN(new_n1553_));
  OAI211_X1 g1188(.A(new_n1553_), .B(new_n554_), .C1(new_n1444_), .C2(new_n1443_), .ZN(new_n1554_));
  AOI21_X1  g1189(.A(new_n1483_), .B1(new_n1492_), .B2(new_n1554_), .ZN(new_n1555_));
  INV_X1    g1190(.A(new_n1485_), .ZN(new_n1556_));
  OAI21_X1  g1191(.A(new_n1552_), .B1(new_n1555_), .B2(new_n1556_), .ZN(new_n1557_));
  INV_X1    g1192(.A(new_n1493_), .ZN(new_n1558_));
  OAI21_X1  g1193(.A(G1497), .B1(new_n1558_), .B2(new_n1452_), .ZN(new_n1559_));
  NAND3_X1  g1194(.A1(new_n1559_), .A2(new_n1485_), .A3(new_n1399_), .ZN(new_n1560_));
  NAND2_X1  g1195(.A1(new_n1557_), .A2(new_n1560_), .ZN(new_n1561_));
  AOI21_X1  g1196(.A(new_n1551_), .B1(new_n1561_), .B2(new_n760_), .ZN(new_n1562_));
  AOI21_X1  g1197(.A(new_n1549_), .B1(new_n1562_), .B2(new_n799_), .ZN(new_n1563_));
  NAND2_X1  g1198(.A1(G94), .A2(G4092), .ZN(new_n1564_));
  INV_X1    g1199(.A(new_n1564_), .ZN(new_n1565_));
  NAND2_X1  g1200(.A1(new_n1368_), .A2(G4091), .ZN(new_n1566_));
  OR2_X1    g1201(.A1(new_n1235_), .A2(G4091), .ZN(new_n1567_));
  XOR2_X1   g1202(.A(new_n1567_), .B(KEYINPUT63), .Z(new_n1568_));
  NAND2_X1  g1203(.A1(new_n1566_), .A2(new_n1568_), .ZN(new_n1569_));
  AOI21_X1  g1204(.A(new_n1565_), .B1(new_n1569_), .B2(new_n755_), .ZN(new_n1570_));
  OAI21_X1  g1205(.A(new_n1563_), .B1(new_n1570_), .B2(new_n983_), .ZN(G767));
  OAI21_X1  g1206(.A(G4090), .B1(G14), .B2(G4089), .ZN(new_n1572_));
  AOI21_X1  g1207(.A(new_n1572_), .B1(new_n1548_), .B2(G4089), .ZN(new_n1573_));
  AOI21_X1  g1208(.A(new_n1573_), .B1(new_n1562_), .B2(new_n843_), .ZN(new_n1574_));
  OAI21_X1  g1209(.A(new_n1574_), .B1(new_n1570_), .B2(new_n1005_), .ZN(G807));
  AOI21_X1  g1210(.A(new_n754_), .B1(new_n1363_), .B2(new_n1367_), .ZN(new_n1576_));
  INV_X1    g1211(.A(new_n1568_), .ZN(new_n1577_));
  OAI21_X1  g1212(.A(new_n755_), .B1(new_n1576_), .B2(new_n1577_), .ZN(new_n1578_));
  AOI21_X1  g1213(.A(new_n1188_), .B1(new_n1578_), .B2(new_n1564_), .ZN(new_n1579_));
  INV_X1    g1214(.A(new_n1551_), .ZN(new_n1580_));
  NAND3_X1  g1215(.A1(new_n1496_), .A2(new_n962_), .A3(new_n1580_), .ZN(new_n1581_));
  INV_X1    g1216(.A(G179), .ZN(new_n1582_));
  NAND2_X1  g1217(.A1(new_n1582_), .A2(G1689), .ZN(new_n1583_));
  OAI211_X1 g1218(.A(new_n1583_), .B(G1690), .C1(G176), .C2(G1689), .ZN(new_n1584_));
  NAND2_X1  g1219(.A1(new_n1581_), .A2(new_n1584_), .ZN(new_n1585_));
  OAI21_X1  g1220(.A(G137), .B1(new_n1579_), .B2(new_n1585_), .ZN(G658));
  AOI21_X1  g1221(.A(new_n1060_), .B1(new_n1578_), .B2(new_n1564_), .ZN(new_n1587_));
  NAND3_X1  g1222(.A1(new_n1496_), .A2(new_n976_), .A3(new_n1580_), .ZN(new_n1588_));
  NAND2_X1  g1223(.A1(new_n1582_), .A2(G1691), .ZN(new_n1589_));
  OAI211_X1 g1224(.A(new_n1589_), .B(G1694), .C1(G176), .C2(G1691), .ZN(new_n1590_));
  NAND2_X1  g1225(.A1(new_n1588_), .A2(new_n1590_), .ZN(new_n1591_));
  OAI21_X1  g1226(.A(G137), .B1(new_n1587_), .B2(new_n1591_), .ZN(G690));
endmodule


