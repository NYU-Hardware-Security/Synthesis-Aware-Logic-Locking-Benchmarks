//Secret key is'0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_c3540" written by ABC on Tue Nov  1 17:40:04 2022

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41,
    G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132,
    G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226,
    G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311,
    G317, G322, G326, G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13,
    G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124,
    G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213,
    G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283,
    G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137_, new_n138_, new_n139_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n980_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1046_, new_n1047_, new_n1048_;
  INV_X1    g000(.A(G58), .ZN(new_n137_));
  INV_X1    g001(.A(G68), .ZN(new_n138_));
  NAND2_X1  g002(.A1(new_n137_), .A2(new_n138_), .ZN(new_n139_));
  NOR3_X1   g003(.A1(new_n139_), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g005(.A1(G1), .A2(G20), .ZN(new_n142_));
  NOR2_X1   g006(.A1(new_n142_), .A2(G13), .ZN(new_n143_));
  INV_X1    g007(.A(new_n143_), .ZN(new_n144_));
  OAI21_X1  g008(.A(G250), .B1(G257), .B2(G264), .ZN(new_n145_));
  NAND2_X1  g009(.A1(new_n139_), .A2(G50), .ZN(new_n146_));
  AND2_X1   g010(.A1(G1), .A2(G13), .ZN(new_n147_));
  NAND2_X1  g011(.A1(new_n147_), .A2(G20), .ZN(new_n148_));
  OAI22_X1  g012(.A1(new_n144_), .A2(new_n145_), .B1(new_n146_), .B2(new_n148_), .ZN(new_n149_));
  AOI22_X1  g013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n150_));
  AOI22_X1  g014(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n151_));
  AOI22_X1  g015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n152_));
  AOI22_X1  g016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n153_));
  NAND4_X1  g017(.A1(new_n150_), .A2(new_n151_), .A3(new_n152_), .A4(new_n153_), .ZN(new_n154_));
  AOI21_X1  g018(.A(new_n149_), .B1(new_n142_), .B2(new_n154_), .ZN(G361));
  XNOR2_X1  g019(.A(G264), .B(G270), .ZN(new_n156_));
  XNOR2_X1  g020(.A(new_n156_), .B(G250), .ZN(new_n157_));
  XNOR2_X1  g021(.A(KEYINPUT0), .B(G257), .ZN(new_n158_));
  XNOR2_X1  g022(.A(new_n157_), .B(new_n158_), .ZN(new_n159_));
  XOR2_X1   g023(.A(G238), .B(G244), .Z(new_n160_));
  XNOR2_X1  g024(.A(G226), .B(G232), .ZN(new_n161_));
  XNOR2_X1  g025(.A(new_n160_), .B(new_n161_), .ZN(new_n162_));
  XNOR2_X1  g026(.A(new_n159_), .B(new_n162_), .ZN(G358));
  XOR2_X1   g027(.A(G87), .B(G97), .Z(new_n164_));
  XNOR2_X1  g028(.A(new_n164_), .B(KEYINPUT1), .ZN(new_n165_));
  XOR2_X1   g029(.A(G107), .B(G116), .Z(new_n166_));
  XNOR2_X1  g030(.A(new_n165_), .B(new_n166_), .ZN(new_n167_));
  XOR2_X1   g031(.A(new_n167_), .B(KEYINPUT2), .Z(new_n168_));
  XNOR2_X1  g032(.A(G68), .B(G77), .ZN(new_n169_));
  XNOR2_X1  g033(.A(G50), .B(G58), .ZN(new_n170_));
  XNOR2_X1  g034(.A(new_n169_), .B(new_n170_), .ZN(new_n171_));
  XNOR2_X1  g035(.A(new_n168_), .B(new_n171_), .ZN(G351));
  NAND2_X1  g036(.A1(G1), .A2(G13), .ZN(new_n173_));
  AOI21_X1  g037(.A(new_n173_), .B1(G33), .B2(G41), .ZN(new_n174_));
  INV_X1    g038(.A(G41), .ZN(new_n175_));
  INV_X1    g039(.A(G45), .ZN(new_n176_));
  AOI21_X1  g040(.A(G1), .B1(new_n175_), .B2(new_n176_), .ZN(new_n177_));
  NOR2_X1   g041(.A1(new_n174_), .A2(new_n177_), .ZN(new_n178_));
  NAND2_X1  g042(.A1(new_n178_), .A2(G226), .ZN(new_n179_));
  NOR2_X1   g043(.A1(G33), .A2(G1698), .ZN(new_n180_));
  NAND2_X1  g044(.A1(new_n180_), .A2(G222), .ZN(new_n181_));
  NAND2_X1  g045(.A1(G33), .A2(G77), .ZN(new_n182_));
  INV_X1    g046(.A(G223), .ZN(new_n183_));
  INV_X1    g047(.A(G33), .ZN(new_n184_));
  NAND2_X1  g048(.A1(new_n184_), .A2(G1698), .ZN(new_n185_));
  OAI211_X1 g049(.A(new_n181_), .B(new_n182_), .C1(new_n183_), .C2(new_n185_), .ZN(new_n186_));
  NAND2_X1  g050(.A1(new_n186_), .A2(new_n174_), .ZN(new_n187_));
  NAND2_X1  g051(.A1(G33), .A2(G41), .ZN(new_n188_));
  NAND3_X1  g052(.A1(new_n188_), .A2(G1), .A3(G13), .ZN(new_n189_));
  AND3_X1   g053(.A1(new_n177_), .A2(new_n189_), .A3(G274), .ZN(new_n190_));
  INV_X1    g054(.A(new_n190_), .ZN(new_n191_));
  NAND3_X1  g055(.A1(new_n179_), .A2(new_n187_), .A3(new_n191_), .ZN(new_n192_));
  INV_X1    g056(.A(G179), .ZN(new_n193_));
  NOR2_X1   g057(.A1(new_n192_), .A2(new_n193_), .ZN(new_n194_));
  AOI21_X1  g058(.A(new_n194_), .B1(G169), .B2(new_n192_), .ZN(new_n195_));
  OAI21_X1  g059(.A(G20), .B1(new_n139_), .B2(G50), .ZN(new_n196_));
  INV_X1    g060(.A(G20), .ZN(new_n197_));
  NAND3_X1  g061(.A1(new_n197_), .A2(new_n184_), .A3(G150), .ZN(new_n198_));
  NAND2_X1  g062(.A1(new_n197_), .A2(G33), .ZN(new_n199_));
  OAI211_X1 g063(.A(new_n196_), .B(new_n198_), .C1(new_n137_), .C2(new_n199_), .ZN(new_n200_));
  NAND3_X1  g064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n201_));
  NAND2_X1  g065(.A1(new_n201_), .A2(new_n173_), .ZN(new_n202_));
  INV_X1    g066(.A(G50), .ZN(new_n203_));
  INV_X1    g067(.A(G1), .ZN(new_n204_));
  NAND2_X1  g068(.A1(new_n204_), .A2(G13), .ZN(new_n205_));
  NOR2_X1   g069(.A1(new_n205_), .A2(new_n197_), .ZN(new_n206_));
  AOI22_X1  g070(.A1(new_n200_), .A2(new_n202_), .B1(new_n203_), .B2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g071(.A1(new_n206_), .A2(new_n202_), .ZN(new_n208_));
  NAND2_X1  g072(.A1(new_n204_), .A2(G20), .ZN(new_n209_));
  NAND3_X1  g073(.A1(new_n208_), .A2(G50), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g074(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g075(.A(new_n211_), .ZN(new_n212_));
  OR2_X1    g076(.A1(new_n195_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g077(.A(KEYINPUT9), .ZN(new_n214_));
  OR2_X1    g078(.A1(new_n192_), .A2(G190), .ZN(new_n215_));
  INV_X1    g079(.A(G200), .ZN(new_n216_));
  NAND2_X1  g080(.A1(new_n192_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g081(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g082(.A(new_n214_), .B1(new_n218_), .B2(new_n212_), .ZN(new_n219_));
  AOI211_X1 g083(.A(KEYINPUT9), .B(new_n211_), .C1(new_n215_), .C2(new_n217_), .ZN(new_n220_));
  OAI21_X1  g084(.A(new_n213_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n222_));
  NAND2_X1  g086(.A1(new_n178_), .A2(G232), .ZN(new_n223_));
  AOI22_X1  g087(.A1(new_n180_), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n224_));
  INV_X1    g088(.A(G1698), .ZN(new_n225_));
  NOR2_X1   g089(.A1(new_n225_), .A2(G33), .ZN(new_n226_));
  NAND2_X1  g090(.A1(new_n226_), .A2(G226), .ZN(new_n227_));
  NAND2_X1  g091(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g092(.A1(new_n228_), .A2(new_n174_), .ZN(new_n229_));
  NAND3_X1  g093(.A1(new_n223_), .A2(new_n229_), .A3(new_n191_), .ZN(new_n230_));
  INV_X1    g094(.A(G190), .ZN(new_n231_));
  OAI21_X1  g095(.A(new_n222_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g096(.A(new_n190_), .B1(G232), .B2(new_n178_), .ZN(new_n233_));
  NAND4_X1  g097(.A1(new_n233_), .A2(KEYINPUT12), .A3(G190), .A4(new_n229_), .ZN(new_n234_));
  NAND2_X1  g098(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g099(.A1(new_n208_), .A2(G58), .A3(new_n209_), .ZN(new_n236_));
  NAND2_X1  g100(.A1(new_n197_), .A2(new_n184_), .ZN(new_n237_));
  INV_X1    g101(.A(G159), .ZN(new_n238_));
  OAI22_X1  g102(.A1(new_n237_), .A2(new_n238_), .B1(new_n199_), .B2(new_n138_), .ZN(new_n239_));
  NAND2_X1  g103(.A1(G58), .A2(G68), .ZN(new_n240_));
  AOI21_X1  g104(.A(new_n197_), .B1(new_n139_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g105(.A(new_n202_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g106(.A(new_n206_), .ZN(new_n243_));
  OAI211_X1 g107(.A(new_n236_), .B(new_n242_), .C1(G58), .C2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g108(.A(new_n244_), .B1(G200), .B2(new_n230_), .ZN(new_n245_));
  NAND2_X1  g109(.A1(new_n235_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g110(.A1(new_n230_), .A2(G169), .ZN(new_n247_));
  OAI21_X1  g111(.A(new_n247_), .B1(new_n193_), .B2(new_n230_), .ZN(new_n248_));
  NAND2_X1  g112(.A1(new_n248_), .A2(new_n244_), .ZN(new_n249_));
  NAND2_X1  g113(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g114(.A1(new_n221_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g115(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g116(.A(new_n190_), .B1(G238), .B2(new_n178_), .ZN(new_n253_));
  NAND2_X1  g117(.A1(new_n180_), .A2(G226), .ZN(new_n254_));
  INV_X1    g118(.A(G97), .ZN(new_n255_));
  INV_X1    g119(.A(G232), .ZN(new_n256_));
  OAI221_X1 g120(.A(new_n254_), .B1(new_n184_), .B2(new_n255_), .C1(new_n256_), .C2(new_n185_), .ZN(new_n257_));
  NAND2_X1  g121(.A1(new_n257_), .A2(new_n174_), .ZN(new_n258_));
  NAND3_X1  g122(.A1(new_n253_), .A2(new_n231_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g123(.A1(new_n178_), .A2(G238), .ZN(new_n260_));
  AND3_X1   g124(.A1(new_n258_), .A2(new_n191_), .A3(new_n260_), .ZN(new_n261_));
  OAI21_X1  g125(.A(new_n259_), .B1(new_n261_), .B2(G200), .ZN(new_n262_));
  OR3_X1    g126(.A1(new_n206_), .A2(KEYINPUT10), .A3(new_n202_), .ZN(new_n263_));
  OAI21_X1  g127(.A(KEYINPUT10), .B1(new_n206_), .B2(new_n202_), .ZN(new_n264_));
  NAND4_X1  g128(.A1(new_n263_), .A2(G68), .A3(new_n264_), .A4(new_n209_), .ZN(new_n265_));
  INV_X1    g129(.A(G13), .ZN(new_n266_));
  AOI211_X1 g130(.A(new_n197_), .B(G68), .C1(new_n201_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g131(.A1(new_n184_), .A2(G50), .ZN(new_n268_));
  AOI21_X1  g132(.A(G20), .B1(new_n268_), .B2(new_n182_), .ZN(new_n269_));
  AOI21_X1  g133(.A(new_n267_), .B1(new_n202_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g134(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g135(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g136(.A1(new_n262_), .A2(new_n272_), .ZN(new_n273_));
  AND3_X1   g137(.A1(new_n253_), .A2(G179), .A3(new_n258_), .ZN(new_n274_));
  INV_X1    g138(.A(G169), .ZN(new_n275_));
  AOI21_X1  g139(.A(new_n275_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n276_));
  OAI21_X1  g140(.A(new_n271_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g141(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g142(.A1(new_n263_), .A2(G77), .A3(new_n264_), .A4(new_n209_), .ZN(new_n279_));
  NAND2_X1  g143(.A1(G20), .A2(G77), .ZN(new_n280_));
  INV_X1    g144(.A(G87), .ZN(new_n281_));
  MUX2_X1   g145(.A(new_n137_), .B(new_n281_), .S(G33), .Z(new_n282_));
  OAI21_X1  g146(.A(new_n280_), .B1(new_n282_), .B2(G20), .ZN(new_n283_));
  INV_X1    g147(.A(G77), .ZN(new_n284_));
  AOI22_X1  g148(.A1(new_n283_), .A2(new_n202_), .B1(new_n284_), .B2(new_n206_), .ZN(new_n285_));
  NAND2_X1  g149(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g150(.A(G244), .ZN(new_n287_));
  NOR3_X1   g151(.A1(new_n174_), .A2(new_n177_), .A3(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g152(.A(new_n288_), .B(KEYINPUT11), .ZN(new_n289_));
  NAND2_X1  g153(.A1(G238), .A2(G1698), .ZN(new_n290_));
  OAI21_X1  g154(.A(new_n290_), .B1(new_n256_), .B2(G1698), .ZN(new_n291_));
  NAND2_X1  g155(.A1(new_n291_), .A2(new_n184_), .ZN(new_n292_));
  INV_X1    g156(.A(G107), .ZN(new_n293_));
  OAI21_X1  g157(.A(new_n292_), .B1(new_n184_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g158(.A(new_n190_), .B1(new_n294_), .B2(new_n174_), .ZN(new_n295_));
  INV_X1    g159(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g160(.A(new_n216_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g161(.A(KEYINPUT11), .ZN(new_n298_));
  XNOR2_X1  g162(.A(new_n288_), .B(new_n298_), .ZN(new_n299_));
  NAND3_X1  g163(.A1(new_n299_), .A2(new_n231_), .A3(new_n295_), .ZN(new_n300_));
  AOI21_X1  g164(.A(new_n286_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g165(.A(new_n301_), .ZN(new_n302_));
  OAI21_X1  g166(.A(G169), .B1(new_n289_), .B2(new_n296_), .ZN(new_n303_));
  NAND3_X1  g167(.A1(new_n299_), .A2(G179), .A3(new_n295_), .ZN(new_n304_));
  NAND2_X1  g168(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g169(.A1(new_n305_), .A2(new_n286_), .ZN(new_n306_));
  NAND2_X1  g170(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g171(.A1(new_n252_), .A2(new_n278_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g172(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g173(.A(KEYINPUT18), .ZN(new_n310_));
  NOR2_X1   g174(.A1(new_n176_), .A2(G1), .ZN(new_n311_));
  NAND4_X1  g175(.A1(new_n189_), .A2(new_n175_), .A3(G274), .A4(new_n311_), .ZN(new_n312_));
  NAND2_X1  g176(.A1(new_n312_), .A2(KEYINPUT5), .ZN(new_n313_));
  INV_X1    g177(.A(G274), .ZN(new_n314_));
  AOI21_X1  g178(.A(new_n314_), .B1(new_n147_), .B2(new_n188_), .ZN(new_n315_));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n316_));
  NAND4_X1  g180(.A1(new_n315_), .A2(new_n316_), .A3(new_n175_), .A4(new_n311_), .ZN(new_n317_));
  NAND2_X1  g181(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g182(.A(KEYINPUT16), .B(G303), .ZN(new_n319_));
  NOR2_X1   g183(.A1(new_n319_), .A2(new_n184_), .ZN(new_n320_));
  NAND2_X1  g184(.A1(new_n225_), .A2(G257), .ZN(new_n321_));
  NAND2_X1  g185(.A1(G264), .A2(G1698), .ZN(new_n322_));
  AOI21_X1  g186(.A(G33), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g187(.A(new_n174_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g188(.A1(new_n204_), .A2(new_n175_), .A3(G45), .ZN(new_n325_));
  AND2_X1   g189(.A1(new_n189_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g190(.A(new_n193_), .B1(new_n326_), .B2(G270), .ZN(new_n327_));
  NAND3_X1  g191(.A1(new_n318_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n329_));
  NAND2_X1  g193(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g194(.A1(new_n318_), .A2(KEYINPUT17), .A3(new_n324_), .A4(new_n327_), .ZN(new_n331_));
  NAND2_X1  g195(.A1(new_n326_), .A2(G270), .ZN(new_n332_));
  NAND3_X1  g196(.A1(new_n318_), .A2(new_n332_), .A3(new_n324_), .ZN(new_n333_));
  AOI22_X1  g197(.A1(new_n330_), .A2(new_n331_), .B1(G169), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g198(.A(G116), .ZN(new_n335_));
  AOI21_X1  g199(.A(new_n335_), .B1(new_n204_), .B2(G33), .ZN(new_n336_));
  NAND3_X1  g200(.A1(new_n263_), .A2(new_n264_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g201(.A(new_n202_), .ZN(new_n338_));
  NOR2_X1   g202(.A1(new_n197_), .A2(G116), .ZN(new_n339_));
  NOR2_X1   g203(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g204(.A(G20), .B1(G33), .B2(G283), .ZN(new_n341_));
  OAI21_X1  g205(.A(new_n341_), .B1(G33), .B2(new_n255_), .ZN(new_n342_));
  INV_X1    g206(.A(new_n205_), .ZN(new_n343_));
  AOI22_X1  g207(.A1(new_n340_), .A2(new_n342_), .B1(new_n343_), .B2(new_n339_), .ZN(new_n344_));
  NAND2_X1  g208(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g209(.A(new_n345_), .ZN(new_n346_));
  OAI21_X1  g210(.A(new_n310_), .B1(new_n334_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g211(.A1(new_n333_), .A2(G169), .ZN(new_n348_));
  INV_X1    g212(.A(G257), .ZN(new_n349_));
  OAI21_X1  g213(.A(new_n322_), .B1(new_n349_), .B2(G1698), .ZN(new_n350_));
  NAND2_X1  g214(.A1(new_n350_), .A2(new_n184_), .ZN(new_n351_));
  OAI21_X1  g215(.A(new_n351_), .B1(new_n184_), .B2(new_n319_), .ZN(new_n352_));
  AOI22_X1  g216(.A1(new_n317_), .A2(new_n313_), .B1(new_n352_), .B2(new_n174_), .ZN(new_n353_));
  AOI21_X1  g217(.A(KEYINPUT17), .B1(new_n353_), .B2(new_n327_), .ZN(new_n354_));
  INV_X1    g218(.A(new_n331_), .ZN(new_n355_));
  OAI21_X1  g219(.A(new_n348_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g220(.A1(new_n356_), .A2(KEYINPUT18), .A3(new_n345_), .ZN(new_n357_));
  NOR2_X1   g221(.A1(new_n333_), .A2(G190), .ZN(new_n358_));
  AOI21_X1  g222(.A(G200), .B1(new_n353_), .B2(new_n332_), .ZN(new_n359_));
  OAI21_X1  g223(.A(new_n346_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AND3_X1   g224(.A1(new_n347_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n361_));
  NAND3_X1  g225(.A1(new_n197_), .A2(G33), .A3(G107), .ZN(new_n362_));
  XOR2_X1   g226(.A(G97), .B(G107), .Z(new_n363_));
  OAI221_X1 g227(.A(new_n362_), .B1(new_n284_), .B2(new_n237_), .C1(new_n363_), .C2(new_n197_), .ZN(new_n364_));
  AOI21_X1  g228(.A(new_n338_), .B1(new_n364_), .B2(KEYINPUT7), .ZN(new_n365_));
  OAI21_X1  g229(.A(new_n365_), .B1(KEYINPUT7), .B2(new_n364_), .ZN(new_n366_));
  OAI21_X1  g230(.A(new_n208_), .B1(G1), .B2(new_n184_), .ZN(new_n367_));
  MUX2_X1   g231(.A(new_n243_), .B(new_n367_), .S(G97), .Z(new_n368_));
  NAND2_X1  g232(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g233(.A1(new_n180_), .A2(G244), .B1(G33), .B2(G283), .ZN(new_n370_));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n371_));
  AOI21_X1  g235(.A(new_n371_), .B1(new_n226_), .B2(G250), .ZN(new_n372_));
  AND4_X1   g236(.A1(new_n371_), .A2(new_n184_), .A3(G250), .A4(G1698), .ZN(new_n373_));
  OAI21_X1  g237(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n375_));
  NAND2_X1  g239(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI211_X1 g240(.A(KEYINPUT4), .B(new_n370_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n377_));
  NAND3_X1  g241(.A1(new_n376_), .A2(new_n174_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g242(.A1(new_n189_), .A2(new_n325_), .A3(G257), .ZN(new_n379_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n380_));
  NAND2_X1  g244(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g245(.A1(new_n189_), .A2(new_n325_), .A3(KEYINPUT6), .A4(G257), .ZN(new_n382_));
  AOI22_X1  g246(.A1(new_n317_), .A2(new_n313_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g247(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g248(.A1(new_n384_), .A2(new_n216_), .ZN(new_n385_));
  NAND3_X1  g249(.A1(new_n378_), .A2(new_n231_), .A3(new_n383_), .ZN(new_n386_));
  AOI21_X1  g250(.A(new_n369_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g251(.A(KEYINPUT8), .ZN(new_n388_));
  NAND2_X1  g252(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g253(.A1(new_n378_), .A2(KEYINPUT8), .A3(new_n383_), .ZN(new_n390_));
  NAND3_X1  g254(.A1(new_n389_), .A2(G179), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g255(.A1(new_n384_), .A2(G169), .ZN(new_n392_));
  NAND2_X1  g256(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g257(.A(new_n387_), .B1(new_n393_), .B2(new_n369_), .ZN(new_n394_));
  NAND3_X1  g258(.A1(new_n343_), .A2(G20), .A3(new_n293_), .ZN(new_n395_));
  NAND2_X1  g259(.A1(new_n335_), .A2(G33), .ZN(new_n396_));
  AOI21_X1  g260(.A(G20), .B1(new_n184_), .B2(new_n281_), .ZN(new_n397_));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n398_));
  OAI21_X1  g262(.A(new_n398_), .B1(new_n197_), .B2(G107), .ZN(new_n399_));
  NAND3_X1  g263(.A1(new_n293_), .A2(KEYINPUT19), .A3(G20), .ZN(new_n400_));
  AOI22_X1  g264(.A1(new_n396_), .A2(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI221_X1 g265(.A(new_n395_), .B1(new_n338_), .B2(new_n401_), .C1(new_n367_), .C2(new_n293_), .ZN(new_n402_));
  INV_X1    g266(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g267(.A(G294), .ZN(new_n404_));
  NOR2_X1   g268(.A1(new_n184_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g269(.A1(G257), .A2(G1698), .ZN(new_n406_));
  INV_X1    g270(.A(G250), .ZN(new_n407_));
  OAI21_X1  g271(.A(new_n406_), .B1(new_n407_), .B2(G1698), .ZN(new_n408_));
  AOI21_X1  g272(.A(new_n405_), .B1(new_n408_), .B2(new_n184_), .ZN(new_n409_));
  INV_X1    g273(.A(new_n409_), .ZN(new_n410_));
  AOI22_X1  g274(.A1(new_n410_), .A2(new_n174_), .B1(G264), .B2(new_n326_), .ZN(new_n411_));
  NAND3_X1  g275(.A1(new_n411_), .A2(G179), .A3(new_n318_), .ZN(new_n412_));
  NAND2_X1  g276(.A1(new_n411_), .A2(new_n318_), .ZN(new_n413_));
  NAND2_X1  g277(.A1(new_n413_), .A2(G169), .ZN(new_n414_));
  AOI21_X1  g278(.A(new_n403_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g279(.A(new_n318_), .ZN(new_n416_));
  NAND2_X1  g280(.A1(new_n326_), .A2(G264), .ZN(new_n417_));
  OAI21_X1  g281(.A(new_n417_), .B1(new_n189_), .B2(new_n409_), .ZN(new_n418_));
  OAI21_X1  g282(.A(new_n216_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g283(.A1(new_n411_), .A2(new_n231_), .A3(new_n318_), .ZN(new_n420_));
  AOI21_X1  g284(.A(new_n402_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g285(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g286(.A1(new_n361_), .A2(new_n394_), .A3(new_n422_), .ZN(new_n423_));
  OAI211_X1 g287(.A(new_n208_), .B(G87), .C1(G1), .C2(new_n184_), .ZN(new_n424_));
  OAI21_X1  g288(.A(new_n424_), .B1(G87), .B2(new_n243_), .ZN(new_n425_));
  NOR2_X1   g289(.A1(new_n237_), .A2(new_n138_), .ZN(new_n426_));
  INV_X1    g290(.A(KEYINPUT13), .ZN(new_n427_));
  NOR3_X1   g291(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n428_));
  AOI21_X1  g292(.A(G20), .B1(G33), .B2(G97), .ZN(new_n429_));
  OAI21_X1  g293(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g294(.A1(new_n197_), .A2(KEYINPUT13), .A3(G33), .A4(G97), .ZN(new_n431_));
  AOI21_X1  g295(.A(new_n426_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g296(.A1(new_n432_), .A2(new_n338_), .ZN(new_n433_));
  NOR2_X1   g297(.A1(new_n425_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n435_));
  NAND3_X1  g299(.A1(new_n189_), .A2(G274), .A3(new_n311_), .ZN(new_n436_));
  NAND2_X1  g300(.A1(new_n204_), .A2(G45), .ZN(new_n437_));
  NAND3_X1  g301(.A1(new_n189_), .A2(G250), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g302(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g303(.A1(new_n225_), .A2(G244), .ZN(new_n440_));
  NOR2_X1   g304(.A1(G238), .A2(G1698), .ZN(new_n441_));
  OAI21_X1  g305(.A(new_n184_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g306(.A1(new_n442_), .A2(KEYINPUT14), .A3(new_n174_), .A4(new_n396_), .ZN(new_n443_));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n444_));
  OR2_X1    g308(.A1(G238), .A2(G1698), .ZN(new_n445_));
  NAND2_X1  g309(.A1(new_n287_), .A2(G1698), .ZN(new_n446_));
  AOI21_X1  g310(.A(G33), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g311(.A1(new_n396_), .A2(new_n147_), .A3(new_n188_), .ZN(new_n448_));
  OAI21_X1  g312(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g313(.A(new_n439_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g314(.A(new_n435_), .B1(new_n450_), .B2(new_n275_), .ZN(new_n451_));
  NAND2_X1  g315(.A1(new_n450_), .A2(G179), .ZN(new_n452_));
  AND2_X1   g316(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g317(.A(new_n450_), .ZN(new_n454_));
  NAND3_X1  g318(.A1(new_n454_), .A2(KEYINPUT15), .A3(G169), .ZN(new_n455_));
  AOI21_X1  g319(.A(new_n434_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  OR2_X1    g320(.A1(new_n425_), .A2(new_n433_), .ZN(new_n457_));
  NAND2_X1  g321(.A1(new_n454_), .A2(new_n216_), .ZN(new_n458_));
  NAND2_X1  g322(.A1(new_n450_), .A2(new_n231_), .ZN(new_n459_));
  AOI21_X1  g323(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NOR4_X1   g324(.A1(new_n309_), .A2(new_n423_), .A3(new_n456_), .A4(new_n460_), .ZN(G372));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n462_));
  OAI21_X1  g326(.A(new_n462_), .B1(new_n252_), .B2(new_n277_), .ZN(new_n463_));
  INV_X1    g327(.A(new_n277_), .ZN(new_n464_));
  NAND3_X1  g328(.A1(new_n251_), .A2(KEYINPUT20), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g329(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g330(.A(new_n286_), .ZN(new_n467_));
  AOI21_X1  g331(.A(new_n467_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n468_));
  NAND4_X1  g332(.A1(new_n468_), .A2(new_n246_), .A3(new_n273_), .A4(new_n277_), .ZN(new_n469_));
  NAND2_X1  g333(.A1(new_n469_), .A2(new_n249_), .ZN(new_n470_));
  OAI21_X1  g334(.A(new_n470_), .B1(new_n220_), .B2(new_n219_), .ZN(new_n471_));
  AND2_X1   g335(.A1(new_n471_), .A2(new_n213_), .ZN(new_n472_));
  NAND2_X1  g336(.A1(new_n466_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g337(.A(new_n473_), .ZN(new_n474_));
  AND3_X1   g338(.A1(new_n378_), .A2(KEYINPUT8), .A3(new_n383_), .ZN(new_n475_));
  AOI21_X1  g339(.A(KEYINPUT8), .B1(new_n378_), .B2(new_n383_), .ZN(new_n476_));
  NOR3_X1   g340(.A1(new_n475_), .A2(new_n476_), .A3(new_n193_), .ZN(new_n477_));
  INV_X1    g341(.A(new_n392_), .ZN(new_n478_));
  OAI21_X1  g342(.A(new_n369_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g343(.A(new_n456_), .ZN(new_n480_));
  NAND2_X1  g344(.A1(new_n330_), .A2(new_n331_), .ZN(new_n481_));
  AOI21_X1  g345(.A(new_n346_), .B1(new_n481_), .B2(new_n348_), .ZN(new_n482_));
  NAND2_X1  g346(.A1(new_n419_), .A2(new_n420_), .ZN(new_n483_));
  NAND2_X1  g347(.A1(new_n483_), .A2(new_n403_), .ZN(new_n484_));
  AOI21_X1  g348(.A(new_n415_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g349(.A(new_n479_), .B(new_n480_), .C1(new_n485_), .C2(new_n387_), .ZN(new_n486_));
  INV_X1    g350(.A(new_n460_), .ZN(new_n487_));
  NAND2_X1  g351(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g352(.A(new_n474_), .B1(new_n309_), .B2(new_n488_), .ZN(G369));
  NAND3_X1  g353(.A1(new_n347_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n490_));
  INV_X1    g354(.A(G213), .ZN(new_n491_));
  NOR3_X1   g355(.A1(new_n205_), .A2(G20), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g356(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g357(.A(G343), .ZN(new_n494_));
  NOR2_X1   g358(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g359(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g360(.A(new_n490_), .B1(new_n346_), .B2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g361(.A1(new_n347_), .A2(new_n357_), .A3(new_n345_), .A4(new_n495_), .ZN(new_n498_));
  NAND2_X1  g362(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g363(.A1(new_n499_), .A2(KEYINPUT21), .ZN(new_n500_));
  NAND2_X1  g364(.A1(new_n402_), .A2(new_n495_), .ZN(new_n501_));
  XNOR2_X1  g365(.A(new_n422_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n503_));
  NAND3_X1  g367(.A1(new_n497_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n504_));
  NAND4_X1  g368(.A1(new_n500_), .A2(G330), .A3(new_n502_), .A4(new_n504_), .ZN(new_n505_));
  NAND2_X1  g369(.A1(new_n347_), .A2(new_n357_), .ZN(new_n506_));
  NAND3_X1  g370(.A1(new_n506_), .A2(new_n422_), .A3(new_n496_), .ZN(new_n507_));
  NAND2_X1  g371(.A1(new_n415_), .A2(new_n496_), .ZN(new_n508_));
  NAND2_X1  g372(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g373(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g374(.A1(new_n505_), .A2(new_n510_), .ZN(G399));
  NOR2_X1   g375(.A1(new_n144_), .A2(G41), .ZN(new_n512_));
  INV_X1    g376(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g377(.A1(new_n428_), .A2(new_n335_), .ZN(new_n514_));
  INV_X1    g378(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g379(.A1(new_n513_), .A2(G1), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g380(.A1(new_n488_), .A2(new_n495_), .ZN(new_n517_));
  INV_X1    g381(.A(G330), .ZN(new_n518_));
  NOR3_X1   g382(.A1(new_n456_), .A2(new_n460_), .A3(new_n495_), .ZN(new_n519_));
  NAND4_X1  g383(.A1(new_n361_), .A2(new_n394_), .A3(new_n519_), .A4(new_n422_), .ZN(new_n520_));
  NOR4_X1   g384(.A1(new_n481_), .A2(new_n413_), .A3(new_n384_), .A4(new_n454_), .ZN(new_n521_));
  NAND4_X1  g385(.A1(new_n413_), .A2(new_n454_), .A3(new_n333_), .A4(new_n193_), .ZN(new_n522_));
  AOI21_X1  g386(.A(new_n522_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n523_));
  OAI21_X1  g387(.A(new_n495_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g388(.A(new_n518_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g389(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  OAI221_X1 g390(.A(new_n516_), .B1(new_n146_), .B2(new_n513_), .C1(new_n526_), .C2(G1), .ZN(G364));
  NOR2_X1   g391(.A1(new_n266_), .A2(G20), .ZN(new_n528_));
  AOI21_X1  g392(.A(new_n204_), .B1(new_n528_), .B2(G45), .ZN(new_n529_));
  INV_X1    g393(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g394(.A1(new_n512_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g395(.A1(new_n143_), .A2(new_n184_), .ZN(new_n532_));
  INV_X1    g396(.A(G355), .ZN(new_n533_));
  OAI22_X1  g397(.A1(new_n532_), .A2(new_n533_), .B1(G116), .B2(new_n143_), .ZN(new_n534_));
  NAND2_X1  g398(.A1(new_n146_), .A2(new_n176_), .ZN(new_n535_));
  OAI21_X1  g399(.A(new_n535_), .B1(new_n171_), .B2(new_n176_), .ZN(new_n536_));
  NOR2_X1   g400(.A1(new_n144_), .A2(new_n184_), .ZN(new_n537_));
  AOI21_X1  g401(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g402(.A1(G13), .A2(G33), .ZN(new_n539_));
  XOR2_X1   g403(.A(new_n539_), .B(KEYINPUT28), .Z(new_n540_));
  NOR2_X1   g404(.A1(new_n540_), .A2(G20), .ZN(new_n541_));
  AOI21_X1  g405(.A(new_n173_), .B1(G20), .B2(new_n275_), .ZN(new_n542_));
  NOR2_X1   g406(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g407(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g408(.A(new_n531_), .B1(new_n538_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g409(.A1(new_n231_), .A2(G20), .ZN(new_n546_));
  OR2_X1    g410(.A1(new_n546_), .A2(KEYINPUT22), .ZN(new_n547_));
  NAND2_X1  g411(.A1(new_n546_), .A2(KEYINPUT22), .ZN(new_n548_));
  NAND2_X1  g412(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NOR3_X1   g413(.A1(new_n197_), .A2(new_n193_), .A3(G200), .ZN(new_n550_));
  NAND2_X1  g414(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NOR4_X1   g415(.A1(new_n197_), .A2(new_n193_), .A3(new_n231_), .A4(new_n216_), .ZN(new_n552_));
  INV_X1    g416(.A(new_n552_), .ZN(new_n553_));
  OAI22_X1  g417(.A1(new_n551_), .A2(new_n137_), .B1(new_n203_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g418(.A(new_n554_), .B(KEYINPUT23), .ZN(new_n555_));
  NOR2_X1   g419(.A1(new_n197_), .A2(new_n231_), .ZN(new_n556_));
  NOR2_X1   g420(.A1(new_n216_), .A2(G179), .ZN(new_n557_));
  NAND2_X1  g421(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g422(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g423(.A1(new_n559_), .A2(G87), .ZN(new_n560_));
  INV_X1    g424(.A(new_n546_), .ZN(new_n561_));
  NAND2_X1  g425(.A1(new_n561_), .A2(new_n557_), .ZN(new_n562_));
  OAI211_X1 g426(.A(new_n560_), .B(new_n184_), .C1(new_n293_), .C2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g427(.A(G20), .B1(G179), .B2(G200), .ZN(new_n564_));
  INV_X1    g428(.A(new_n564_), .ZN(new_n565_));
  NOR2_X1   g429(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g430(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g431(.A1(new_n550_), .A2(new_n231_), .ZN(new_n568_));
  OAI22_X1  g432(.A1(new_n567_), .A2(new_n255_), .B1(new_n284_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g433(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g434(.A1(new_n549_), .A2(new_n565_), .ZN(new_n571_));
  NOR3_X1   g435(.A1(new_n197_), .A2(new_n193_), .A3(new_n216_), .ZN(new_n572_));
  NAND3_X1  g436(.A1(new_n547_), .A2(new_n572_), .A3(new_n548_), .ZN(new_n573_));
  INV_X1    g437(.A(new_n573_), .ZN(new_n574_));
  AOI22_X1  g438(.A1(new_n571_), .A2(G159), .B1(new_n574_), .B2(G68), .ZN(new_n575_));
  NAND3_X1  g439(.A1(new_n555_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g440(.A(G283), .ZN(new_n577_));
  NOR2_X1   g441(.A1(new_n562_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g442(.A(new_n578_), .B(KEYINPUT25), .ZN(new_n579_));
  NAND2_X1  g443(.A1(new_n552_), .A2(G326), .ZN(new_n580_));
  INV_X1    g444(.A(G311), .ZN(new_n581_));
  OAI221_X1 g445(.A(new_n580_), .B1(new_n581_), .B2(new_n568_), .C1(new_n319_), .C2(new_n558_), .ZN(new_n582_));
  INV_X1    g446(.A(G322), .ZN(new_n583_));
  INV_X1    g447(.A(G317), .ZN(new_n584_));
  OAI22_X1  g448(.A1(new_n551_), .A2(new_n583_), .B1(new_n584_), .B2(new_n573_), .ZN(new_n585_));
  AOI211_X1 g449(.A(new_n582_), .B(new_n585_), .C1(G294), .C2(new_n566_), .ZN(new_n586_));
  XNOR2_X1  g450(.A(new_n586_), .B(KEYINPUT24), .ZN(new_n587_));
  AOI211_X1 g451(.A(new_n579_), .B(new_n587_), .C1(G329), .C2(new_n571_), .ZN(new_n588_));
  INV_X1    g452(.A(KEYINPUT26), .ZN(new_n589_));
  AND2_X1   g453(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g454(.A(G33), .B1(new_n588_), .B2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g455(.A(new_n576_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g456(.A1(new_n592_), .A2(KEYINPUT27), .ZN(new_n593_));
  INV_X1    g457(.A(new_n542_), .ZN(new_n594_));
  AOI21_X1  g458(.A(new_n594_), .B1(new_n592_), .B2(KEYINPUT27), .ZN(new_n595_));
  AOI21_X1  g459(.A(new_n545_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  AND2_X1   g460(.A1(new_n500_), .A2(new_n504_), .ZN(new_n597_));
  INV_X1    g461(.A(new_n541_), .ZN(new_n598_));
  OR2_X1    g462(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OR2_X1    g463(.A1(new_n597_), .A2(G330), .ZN(new_n600_));
  NAND3_X1  g464(.A1(new_n500_), .A2(G330), .A3(new_n504_), .ZN(new_n601_));
  INV_X1    g465(.A(new_n531_), .ZN(new_n602_));
  AND2_X1   g466(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI22_X1  g467(.A1(new_n596_), .A2(new_n599_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g468(.A(new_n604_), .ZN(G396));
  NOR2_X1   g469(.A1(new_n307_), .A2(new_n495_), .ZN(new_n606_));
  NAND2_X1  g470(.A1(new_n479_), .A2(new_n480_), .ZN(new_n607_));
  NAND3_X1  g471(.A1(new_n484_), .A2(new_n356_), .A3(new_n345_), .ZN(new_n608_));
  INV_X1    g472(.A(new_n415_), .ZN(new_n609_));
  AOI21_X1  g473(.A(new_n387_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI211_X1 g474(.A(new_n487_), .B(new_n606_), .C1(new_n607_), .C2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g475(.A1(new_n286_), .A2(new_n495_), .ZN(new_n612_));
  OAI21_X1  g476(.A(new_n612_), .B1(new_n301_), .B2(new_n468_), .ZN(new_n613_));
  OAI21_X1  g477(.A(new_n613_), .B1(new_n468_), .B2(new_n612_), .ZN(new_n614_));
  INV_X1    g478(.A(new_n614_), .ZN(new_n615_));
  OAI21_X1  g479(.A(new_n611_), .B1(new_n517_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g480(.A(new_n616_), .B(KEYINPUT29), .ZN(new_n617_));
  AOI21_X1  g481(.A(new_n531_), .B1(new_n617_), .B2(new_n525_), .ZN(new_n618_));
  OAI21_X1  g482(.A(new_n618_), .B1(new_n525_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g483(.A1(new_n542_), .A2(new_n539_), .ZN(new_n620_));
  AOI21_X1  g484(.A(new_n602_), .B1(new_n284_), .B2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g485(.A1(new_n562_), .A2(new_n281_), .ZN(new_n622_));
  INV_X1    g486(.A(G303), .ZN(new_n623_));
  OAI21_X1  g487(.A(G33), .B1(new_n553_), .B2(new_n623_), .ZN(new_n624_));
  AOI211_X1 g488(.A(new_n622_), .B(new_n624_), .C1(G107), .C2(new_n559_), .ZN(new_n625_));
  INV_X1    g489(.A(new_n568_), .ZN(new_n626_));
  AOI22_X1  g490(.A1(new_n626_), .A2(G116), .B1(G97), .B2(new_n566_), .ZN(new_n627_));
  INV_X1    g491(.A(new_n551_), .ZN(new_n628_));
  NAND2_X1  g492(.A1(new_n628_), .A2(G294), .ZN(new_n629_));
  AOI22_X1  g493(.A1(new_n571_), .A2(G311), .B1(new_n574_), .B2(G283), .ZN(new_n630_));
  NAND4_X1  g494(.A1(new_n625_), .A2(new_n627_), .A3(new_n629_), .A4(new_n630_), .ZN(new_n631_));
  INV_X1    g495(.A(G143), .ZN(new_n632_));
  INV_X1    g496(.A(G150), .ZN(new_n633_));
  OAI22_X1  g497(.A1(new_n551_), .A2(new_n632_), .B1(new_n633_), .B2(new_n573_), .ZN(new_n634_));
  AOI21_X1  g498(.A(new_n634_), .B1(G132), .B2(new_n571_), .ZN(new_n635_));
  AOI21_X1  g499(.A(G33), .B1(new_n552_), .B2(G137), .ZN(new_n636_));
  INV_X1    g500(.A(new_n562_), .ZN(new_n637_));
  AOI22_X1  g501(.A1(new_n637_), .A2(G68), .B1(new_n559_), .B2(G50), .ZN(new_n638_));
  AOI22_X1  g502(.A1(new_n626_), .A2(G159), .B1(G58), .B2(new_n566_), .ZN(new_n639_));
  NAND4_X1  g503(.A1(new_n635_), .A2(new_n636_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n640_));
  NAND2_X1  g504(.A1(new_n631_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g505(.A1(new_n641_), .A2(KEYINPUT30), .ZN(new_n642_));
  NAND2_X1  g506(.A1(new_n642_), .A2(new_n542_), .ZN(new_n643_));
  NOR2_X1   g507(.A1(new_n641_), .A2(KEYINPUT30), .ZN(new_n644_));
  OAI221_X1 g508(.A(new_n621_), .B1(new_n643_), .B2(new_n644_), .C1(new_n615_), .C2(new_n540_), .ZN(new_n645_));
  NAND2_X1  g509(.A1(new_n619_), .A2(new_n645_), .ZN(G384));
  NOR2_X1   g510(.A1(new_n528_), .A2(new_n204_), .ZN(new_n647_));
  AOI21_X1  g511(.A(new_n473_), .B1(new_n308_), .B2(new_n517_), .ZN(new_n648_));
  NAND2_X1  g512(.A1(new_n271_), .A2(new_n495_), .ZN(new_n649_));
  NAND3_X1  g513(.A1(new_n273_), .A2(new_n277_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g514(.A(KEYINPUT32), .ZN(new_n651_));
  NAND2_X1  g515(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g516(.A1(new_n273_), .A2(KEYINPUT32), .A3(new_n277_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g517(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OR3_X1    g518(.A1(new_n277_), .A2(KEYINPUT31), .A3(new_n496_), .ZN(new_n655_));
  OAI21_X1  g519(.A(KEYINPUT31), .B1(new_n277_), .B2(new_n496_), .ZN(new_n656_));
  NAND2_X1  g520(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g521(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g522(.A1(new_n250_), .A2(new_n244_), .A3(new_n492_), .ZN(new_n659_));
  NAND2_X1  g523(.A1(new_n244_), .A2(new_n492_), .ZN(new_n660_));
  NAND3_X1  g524(.A1(new_n246_), .A2(new_n249_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g525(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g526(.A1(new_n306_), .A2(new_n495_), .ZN(new_n663_));
  NAND3_X1  g527(.A1(new_n658_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NOR2_X1   g528(.A1(new_n249_), .A2(new_n492_), .ZN(new_n665_));
  NOR2_X1   g529(.A1(new_n277_), .A2(new_n495_), .ZN(new_n666_));
  AOI21_X1  g530(.A(new_n665_), .B1(new_n662_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g531(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  AOI22_X1  g532(.A1(new_n652_), .A2(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n669_));
  NAND4_X1  g533(.A1(new_n486_), .A2(new_n487_), .A3(new_n606_), .A4(new_n662_), .ZN(new_n670_));
  AOI21_X1  g534(.A(new_n669_), .B1(new_n670_), .B2(KEYINPUT33), .ZN(new_n671_));
  INV_X1    g535(.A(new_n387_), .ZN(new_n672_));
  NOR3_X1   g536(.A1(new_n334_), .A2(new_n421_), .A3(new_n346_), .ZN(new_n673_));
  OAI21_X1  g537(.A(new_n672_), .B1(new_n673_), .B2(new_n415_), .ZN(new_n674_));
  AOI21_X1  g538(.A(new_n456_), .B1(new_n393_), .B2(new_n369_), .ZN(new_n675_));
  AOI21_X1  g539(.A(new_n460_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g540(.A(KEYINPUT33), .ZN(new_n677_));
  NAND4_X1  g541(.A1(new_n676_), .A2(new_n677_), .A3(new_n606_), .A4(new_n662_), .ZN(new_n678_));
  AOI21_X1  g542(.A(new_n668_), .B1(new_n671_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g543(.A(new_n648_), .B(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g544(.A(new_n250_), .B(new_n660_), .ZN(new_n681_));
  NOR3_X1   g545(.A1(new_n669_), .A2(new_n681_), .A3(new_n614_), .ZN(new_n682_));
  XOR2_X1   g546(.A(new_n308_), .B(new_n682_), .Z(new_n683_));
  NAND2_X1  g547(.A1(new_n683_), .A2(new_n525_), .ZN(new_n684_));
  AOI21_X1  g548(.A(new_n647_), .B1(new_n680_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g549(.A(new_n685_), .B1(new_n680_), .B2(new_n684_), .ZN(new_n686_));
  NAND2_X1  g550(.A1(new_n240_), .A2(G77), .ZN(new_n687_));
  OAI22_X1  g551(.A1(new_n146_), .A2(new_n687_), .B1(G50), .B2(new_n138_), .ZN(new_n688_));
  NOR2_X1   g552(.A1(new_n204_), .A2(G13), .ZN(new_n689_));
  NOR2_X1   g553(.A1(new_n148_), .A2(new_n335_), .ZN(new_n690_));
  AOI22_X1  g554(.A1(new_n688_), .A2(new_n689_), .B1(new_n363_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g555(.A1(new_n686_), .A2(new_n691_), .ZN(G367));
  NAND3_X1  g556(.A1(new_n393_), .A2(new_n369_), .A3(new_n496_), .ZN(new_n693_));
  NAND2_X1  g557(.A1(new_n369_), .A2(new_n495_), .ZN(new_n694_));
  INV_X1    g558(.A(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g559(.A(new_n394_), .B(new_n695_), .ZN(new_n696_));
  OAI21_X1  g560(.A(new_n693_), .B1(new_n696_), .B2(new_n510_), .ZN(new_n697_));
  NAND2_X1  g561(.A1(new_n697_), .A2(KEYINPUT34), .ZN(new_n698_));
  NOR2_X1   g562(.A1(new_n456_), .A2(new_n460_), .ZN(new_n699_));
  NAND2_X1  g563(.A1(new_n457_), .A2(new_n495_), .ZN(new_n700_));
  XNOR2_X1  g564(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  INV_X1    g565(.A(KEYINPUT34), .ZN(new_n702_));
  OAI211_X1 g566(.A(new_n702_), .B(new_n693_), .C1(new_n696_), .C2(new_n510_), .ZN(new_n703_));
  NAND3_X1  g567(.A1(new_n698_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  OR3_X1    g568(.A1(new_n697_), .A2(KEYINPUT34), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g569(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g570(.A(new_n505_), .ZN(new_n707_));
  NAND2_X1  g571(.A1(new_n479_), .A2(new_n672_), .ZN(new_n708_));
  NAND2_X1  g572(.A1(new_n708_), .A2(new_n695_), .ZN(new_n709_));
  NAND2_X1  g573(.A1(new_n394_), .A2(new_n694_), .ZN(new_n710_));
  NAND2_X1  g574(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g575(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g576(.A(new_n706_), .B(new_n712_), .ZN(new_n713_));
  INV_X1    g577(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g578(.A1(new_n711_), .A2(KEYINPUT35), .ZN(new_n715_));
  INV_X1    g579(.A(KEYINPUT35), .ZN(new_n716_));
  NAND3_X1  g580(.A1(new_n709_), .A2(new_n716_), .A3(new_n710_), .ZN(new_n717_));
  NAND3_X1  g581(.A1(new_n715_), .A2(new_n717_), .A3(new_n509_), .ZN(new_n718_));
  NAND3_X1  g582(.A1(new_n696_), .A2(new_n510_), .A3(new_n716_), .ZN(new_n719_));
  NAND2_X1  g583(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g584(.A1(new_n720_), .A2(new_n707_), .ZN(new_n721_));
  NAND3_X1  g585(.A1(new_n718_), .A2(new_n505_), .A3(new_n719_), .ZN(new_n722_));
  AND2_X1   g586(.A1(new_n347_), .A2(new_n357_), .ZN(new_n723_));
  NOR2_X1   g587(.A1(new_n723_), .A2(new_n495_), .ZN(new_n724_));
  OAI21_X1  g588(.A(new_n507_), .B1(new_n502_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g589(.A(new_n725_), .ZN(new_n726_));
  NAND2_X1  g590(.A1(new_n601_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g591(.A1(new_n597_), .A2(G330), .A3(new_n725_), .ZN(new_n728_));
  AOI22_X1  g592(.A1(new_n721_), .A2(new_n722_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  OR2_X1    g593(.A1(new_n517_), .A2(new_n525_), .ZN(new_n730_));
  OAI21_X1  g594(.A(new_n512_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g595(.A1(new_n731_), .A2(new_n529_), .ZN(new_n732_));
  NAND2_X1  g596(.A1(new_n714_), .A2(new_n732_), .ZN(new_n733_));
  OR2_X1    g597(.A1(new_n701_), .A2(new_n598_), .ZN(new_n734_));
  NOR3_X1   g598(.A1(new_n159_), .A2(new_n184_), .A3(new_n144_), .ZN(new_n735_));
  OAI21_X1  g599(.A(new_n543_), .B1(new_n281_), .B2(new_n143_), .ZN(new_n736_));
  OAI21_X1  g600(.A(new_n531_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AOI22_X1  g601(.A1(new_n571_), .A2(G137), .B1(new_n574_), .B2(G159), .ZN(new_n738_));
  OAI21_X1  g602(.A(new_n738_), .B1(new_n633_), .B2(new_n551_), .ZN(new_n739_));
  OAI21_X1  g603(.A(new_n184_), .B1(new_n558_), .B2(new_n137_), .ZN(new_n740_));
  NAND2_X1  g604(.A1(new_n637_), .A2(G77), .ZN(new_n741_));
  OAI21_X1  g605(.A(new_n741_), .B1(new_n553_), .B2(new_n632_), .ZN(new_n742_));
  NAND2_X1  g606(.A1(new_n566_), .A2(G68), .ZN(new_n743_));
  OAI21_X1  g607(.A(new_n743_), .B1(new_n203_), .B2(new_n568_), .ZN(new_n744_));
  NOR4_X1   g608(.A1(new_n739_), .A2(new_n740_), .A3(new_n742_), .A4(new_n744_), .ZN(new_n745_));
  OR2_X1    g609(.A1(new_n745_), .A2(KEYINPUT36), .ZN(new_n746_));
  NAND2_X1  g610(.A1(new_n745_), .A2(KEYINPUT36), .ZN(new_n747_));
  OAI22_X1  g611(.A1(new_n567_), .A2(new_n293_), .B1(new_n577_), .B2(new_n568_), .ZN(new_n748_));
  OAI21_X1  g612(.A(G33), .B1(new_n553_), .B2(new_n581_), .ZN(new_n749_));
  OAI22_X1  g613(.A1(new_n562_), .A2(new_n255_), .B1(new_n558_), .B2(new_n335_), .ZN(new_n750_));
  NOR3_X1   g614(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g615(.A(KEYINPUT37), .B(G294), .ZN(new_n752_));
  INV_X1    g616(.A(new_n752_), .ZN(new_n753_));
  AOI22_X1  g617(.A1(new_n571_), .A2(G317), .B1(new_n574_), .B2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g618(.A(new_n751_), .B(new_n754_), .C1(new_n623_), .C2(new_n551_), .ZN(new_n755_));
  NAND3_X1  g619(.A1(new_n746_), .A2(new_n747_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g620(.A(new_n737_), .B1(new_n756_), .B2(new_n542_), .ZN(new_n757_));
  NAND2_X1  g621(.A1(new_n734_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g622(.A1(new_n733_), .A2(new_n758_), .ZN(G387));
  AOI21_X1  g623(.A(new_n730_), .B1(new_n728_), .B2(new_n727_), .ZN(new_n760_));
  NOR2_X1   g624(.A1(new_n760_), .A2(new_n513_), .ZN(new_n761_));
  NAND2_X1  g625(.A1(new_n728_), .A2(new_n727_), .ZN(new_n762_));
  OAI21_X1  g626(.A(new_n761_), .B1(new_n526_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g627(.A1(new_n762_), .A2(new_n530_), .ZN(new_n764_));
  AOI21_X1  g628(.A(G45), .B1(G68), .B2(G77), .ZN(new_n765_));
  NAND3_X1  g629(.A1(new_n765_), .A2(new_n203_), .A3(G58), .ZN(new_n766_));
  OAI221_X1 g630(.A(new_n537_), .B1(new_n514_), .B2(new_n766_), .C1(new_n162_), .C2(new_n176_), .ZN(new_n767_));
  XOR2_X1   g631(.A(new_n767_), .B(KEYINPUT40), .Z(new_n768_));
  OAI221_X1 g632(.A(new_n768_), .B1(G107), .B2(new_n143_), .C1(new_n515_), .C2(new_n532_), .ZN(new_n769_));
  AOI21_X1  g633(.A(new_n602_), .B1(new_n769_), .B2(new_n543_), .ZN(new_n770_));
  NAND2_X1  g634(.A1(new_n571_), .A2(G326), .ZN(new_n771_));
  XOR2_X1   g635(.A(new_n771_), .B(KEYINPUT39), .Z(new_n772_));
  OAI22_X1  g636(.A1(new_n567_), .A2(new_n577_), .B1(new_n319_), .B2(new_n568_), .ZN(new_n773_));
  OAI22_X1  g637(.A1(new_n553_), .A2(new_n583_), .B1(new_n558_), .B2(new_n752_), .ZN(new_n774_));
  OAI21_X1  g638(.A(G33), .B1(new_n562_), .B2(new_n335_), .ZN(new_n775_));
  NOR3_X1   g639(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AOI22_X1  g640(.A1(new_n628_), .A2(G317), .B1(G311), .B2(new_n574_), .ZN(new_n777_));
  NAND3_X1  g641(.A1(new_n772_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g642(.A(new_n184_), .B1(new_n562_), .B2(new_n255_), .ZN(new_n779_));
  OAI22_X1  g643(.A1(new_n567_), .A2(new_n281_), .B1(new_n138_), .B2(new_n568_), .ZN(new_n780_));
  AOI211_X1 g644(.A(new_n779_), .B(new_n780_), .C1(G77), .C2(new_n559_), .ZN(new_n781_));
  OAI22_X1  g645(.A1(new_n551_), .A2(new_n203_), .B1(new_n238_), .B2(new_n553_), .ZN(new_n782_));
  OR2_X1    g646(.A1(new_n782_), .A2(KEYINPUT38), .ZN(new_n783_));
  NAND2_X1  g647(.A1(new_n782_), .A2(KEYINPUT38), .ZN(new_n784_));
  AOI22_X1  g648(.A1(new_n571_), .A2(G150), .B1(new_n574_), .B2(G58), .ZN(new_n785_));
  NAND4_X1  g649(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .A4(new_n785_), .ZN(new_n786_));
  AND2_X1   g650(.A1(new_n778_), .A2(new_n786_), .ZN(new_n787_));
  OAI221_X1 g651(.A(new_n770_), .B1(new_n502_), .B2(new_n598_), .C1(new_n594_), .C2(new_n787_), .ZN(new_n788_));
  AND2_X1   g652(.A1(new_n764_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g653(.A1(new_n763_), .A2(new_n789_), .ZN(G393));
  AOI21_X1  g654(.A(new_n529_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n791_));
  INV_X1    g655(.A(KEYINPUT43), .ZN(new_n792_));
  AND2_X1   g656(.A1(new_n167_), .A2(new_n537_), .ZN(new_n793_));
  OAI21_X1  g657(.A(new_n543_), .B1(new_n255_), .B2(new_n143_), .ZN(new_n794_));
  OAI21_X1  g658(.A(new_n531_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI22_X1  g659(.A1(new_n567_), .A2(new_n284_), .B1(new_n137_), .B2(new_n568_), .ZN(new_n796_));
  OAI22_X1  g660(.A1(new_n553_), .A2(new_n633_), .B1(new_n558_), .B2(new_n138_), .ZN(new_n797_));
  NOR4_X1   g661(.A1(new_n796_), .A2(new_n797_), .A3(G33), .A4(new_n622_), .ZN(new_n798_));
  AOI22_X1  g662(.A1(new_n628_), .A2(G159), .B1(new_n571_), .B2(G143), .ZN(new_n799_));
  OAI211_X1 g663(.A(new_n798_), .B(new_n799_), .C1(new_n203_), .C2(new_n573_), .ZN(new_n800_));
  NOR2_X1   g664(.A1(new_n567_), .A2(new_n335_), .ZN(new_n801_));
  OAI22_X1  g665(.A1(new_n553_), .A2(new_n584_), .B1(new_n558_), .B2(new_n577_), .ZN(new_n802_));
  AOI211_X1 g666(.A(new_n801_), .B(new_n802_), .C1(new_n626_), .C2(new_n753_), .ZN(new_n803_));
  OAI221_X1 g667(.A(new_n803_), .B1(new_n581_), .B2(new_n551_), .C1(new_n319_), .C2(new_n573_), .ZN(new_n804_));
  INV_X1    g668(.A(KEYINPUT42), .ZN(new_n805_));
  NAND2_X1  g669(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g670(.A(G33), .B1(new_n562_), .B2(new_n293_), .ZN(new_n807_));
  AOI21_X1  g671(.A(new_n807_), .B1(new_n571_), .B2(G322), .ZN(new_n808_));
  NAND2_X1  g672(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g673(.A1(new_n804_), .A2(new_n805_), .ZN(new_n810_));
  OAI21_X1  g674(.A(new_n800_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g675(.A(new_n795_), .B1(new_n811_), .B2(new_n542_), .ZN(new_n812_));
  OAI21_X1  g676(.A(new_n812_), .B1(new_n711_), .B2(new_n598_), .ZN(new_n813_));
  INV_X1    g677(.A(new_n813_), .ZN(new_n814_));
  OR3_X1    g678(.A1(new_n791_), .A2(new_n792_), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g679(.A(new_n792_), .B1(new_n791_), .B2(new_n814_), .ZN(new_n816_));
  NAND2_X1  g680(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g681(.A1(new_n721_), .A2(new_n722_), .ZN(new_n818_));
  INV_X1    g682(.A(KEYINPUT41), .ZN(new_n819_));
  AOI21_X1  g683(.A(new_n819_), .B1(new_n720_), .B2(new_n707_), .ZN(new_n820_));
  OR3_X1    g684(.A1(new_n818_), .A2(new_n760_), .A3(new_n820_), .ZN(new_n821_));
  OAI21_X1  g685(.A(new_n818_), .B1(new_n760_), .B2(new_n820_), .ZN(new_n822_));
  NAND3_X1  g686(.A1(new_n821_), .A2(new_n512_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g687(.A1(new_n817_), .A2(new_n823_), .ZN(G390));
  INV_X1    g688(.A(new_n620_), .ZN(new_n825_));
  OAI21_X1  g689(.A(new_n531_), .B1(G58), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g690(.A1(new_n681_), .A2(new_n539_), .ZN(new_n827_));
  XOR2_X1   g691(.A(new_n827_), .B(KEYINPUT49), .Z(new_n828_));
  AOI22_X1  g692(.A1(new_n571_), .A2(G294), .B1(new_n574_), .B2(G107), .ZN(new_n829_));
  OAI21_X1  g693(.A(new_n829_), .B1(new_n335_), .B2(new_n551_), .ZN(new_n830_));
  AOI22_X1  g694(.A1(new_n626_), .A2(G97), .B1(G77), .B2(new_n566_), .ZN(new_n831_));
  AOI22_X1  g695(.A1(new_n637_), .A2(G68), .B1(new_n552_), .B2(G283), .ZN(new_n832_));
  NAND4_X1  g696(.A1(new_n831_), .A2(new_n832_), .A3(G33), .A4(new_n560_), .ZN(new_n833_));
  AOI22_X1  g697(.A1(new_n571_), .A2(G125), .B1(new_n574_), .B2(G137), .ZN(new_n834_));
  NOR2_X1   g698(.A1(new_n562_), .A2(new_n203_), .ZN(new_n835_));
  XNOR2_X1  g699(.A(new_n835_), .B(KEYINPUT48), .ZN(new_n836_));
  NAND2_X1  g700(.A1(new_n628_), .A2(G132), .ZN(new_n837_));
  NAND3_X1  g701(.A1(new_n834_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI22_X1  g702(.A1(new_n626_), .A2(G143), .B1(G159), .B2(new_n566_), .ZN(new_n839_));
  AOI21_X1  g703(.A(G33), .B1(new_n552_), .B2(G128), .ZN(new_n840_));
  OAI211_X1 g704(.A(new_n839_), .B(new_n840_), .C1(new_n633_), .C2(new_n558_), .ZN(new_n841_));
  OAI22_X1  g705(.A1(new_n830_), .A2(new_n833_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n842_));
  AOI211_X1 g706(.A(new_n826_), .B(new_n828_), .C1(new_n542_), .C2(new_n842_), .ZN(new_n843_));
  AOI211_X1 g707(.A(new_n518_), .B(new_n614_), .C1(new_n520_), .C2(new_n524_), .ZN(new_n844_));
  INV_X1    g708(.A(new_n663_), .ZN(new_n845_));
  NAND2_X1  g709(.A1(new_n611_), .A2(new_n845_), .ZN(new_n846_));
  OAI22_X1  g710(.A1(new_n662_), .A2(KEYINPUT45), .B1(new_n277_), .B2(new_n495_), .ZN(new_n847_));
  OAI211_X1 g711(.A(new_n844_), .B(new_n658_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g712(.A(new_n847_), .B1(new_n846_), .B2(new_n658_), .ZN(new_n849_));
  NAND2_X1  g713(.A1(new_n520_), .A2(new_n524_), .ZN(new_n850_));
  NAND4_X1  g714(.A1(new_n850_), .A2(G330), .A3(new_n615_), .A4(new_n658_), .ZN(new_n851_));
  NAND2_X1  g715(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g716(.A1(new_n681_), .A2(KEYINPUT44), .ZN(new_n853_));
  AND2_X1   g717(.A1(new_n853_), .A2(KEYINPUT45), .ZN(new_n854_));
  AND3_X1   g718(.A1(new_n848_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g719(.A(new_n854_), .B1(new_n848_), .B2(new_n852_), .ZN(new_n856_));
  NOR2_X1   g720(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g721(.A(new_n843_), .B1(new_n857_), .B2(new_n530_), .ZN(new_n858_));
  INV_X1    g722(.A(new_n854_), .ZN(new_n859_));
  AND2_X1   g723(.A1(new_n849_), .A2(new_n851_), .ZN(new_n860_));
  NOR2_X1   g724(.A1(new_n849_), .A2(new_n851_), .ZN(new_n861_));
  OAI21_X1  g725(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g726(.A1(new_n848_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n863_));
  NAND2_X1  g727(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g728(.A(new_n473_), .B1(new_n308_), .B2(new_n730_), .ZN(new_n865_));
  NAND3_X1  g729(.A1(new_n611_), .A2(new_n658_), .A3(new_n845_), .ZN(new_n866_));
  INV_X1    g730(.A(KEYINPUT47), .ZN(new_n867_));
  NAND2_X1  g731(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g732(.A1(new_n846_), .A2(new_n669_), .ZN(new_n869_));
  NAND2_X1  g733(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI211_X1 g734(.A(KEYINPUT47), .B(new_n658_), .C1(new_n611_), .C2(new_n845_), .ZN(new_n871_));
  INV_X1    g735(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g736(.A(new_n844_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g737(.A1(new_n866_), .A2(new_n525_), .A3(new_n615_), .ZN(new_n874_));
  AOI21_X1  g738(.A(KEYINPUT46), .B1(new_n846_), .B2(new_n669_), .ZN(new_n875_));
  INV_X1    g739(.A(KEYINPUT46), .ZN(new_n876_));
  AOI211_X1 g740(.A(new_n876_), .B(new_n658_), .C1(new_n611_), .C2(new_n845_), .ZN(new_n877_));
  NOR3_X1   g741(.A1(new_n874_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g742(.A(new_n865_), .B1(new_n873_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g743(.A(new_n512_), .B1(new_n864_), .B2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g744(.A(new_n663_), .B1(new_n676_), .B2(new_n606_), .ZN(new_n881_));
  OAI21_X1  g745(.A(new_n876_), .B1(new_n881_), .B2(new_n658_), .ZN(new_n882_));
  NAND3_X1  g746(.A1(new_n846_), .A2(KEYINPUT46), .A3(new_n669_), .ZN(new_n883_));
  NAND4_X1  g747(.A1(new_n882_), .A2(new_n844_), .A3(new_n883_), .A4(new_n866_), .ZN(new_n884_));
  AOI21_X1  g748(.A(new_n871_), .B1(new_n869_), .B2(new_n868_), .ZN(new_n885_));
  OAI21_X1  g749(.A(new_n884_), .B1(new_n885_), .B2(new_n844_), .ZN(new_n886_));
  AOI22_X1  g750(.A1(new_n886_), .A2(new_n865_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n887_));
  OAI21_X1  g751(.A(new_n858_), .B1(new_n880_), .B2(new_n887_), .ZN(G378));
  NAND2_X1  g752(.A1(new_n211_), .A2(new_n492_), .ZN(new_n889_));
  INV_X1    g753(.A(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g754(.A(new_n221_), .B(new_n890_), .ZN(new_n891_));
  NOR2_X1   g755(.A1(new_n891_), .A2(new_n540_), .ZN(new_n892_));
  AOI22_X1  g756(.A1(new_n571_), .A2(G283), .B1(new_n574_), .B2(G97), .ZN(new_n893_));
  OAI21_X1  g757(.A(new_n893_), .B1(new_n293_), .B2(new_n551_), .ZN(new_n894_));
  OAI211_X1 g758(.A(G33), .B(new_n175_), .C1(new_n558_), .C2(new_n284_), .ZN(new_n895_));
  NAND2_X1  g759(.A1(new_n637_), .A2(G58), .ZN(new_n896_));
  OAI21_X1  g760(.A(new_n896_), .B1(new_n553_), .B2(new_n335_), .ZN(new_n897_));
  OAI21_X1  g761(.A(new_n743_), .B1(new_n281_), .B2(new_n568_), .ZN(new_n898_));
  NOR4_X1   g762(.A1(new_n894_), .A2(new_n895_), .A3(new_n897_), .A4(new_n898_), .ZN(new_n899_));
  XOR2_X1   g763(.A(new_n899_), .B(KEYINPUT53), .Z(new_n900_));
  AOI211_X1 g764(.A(G33), .B(G41), .C1(new_n559_), .C2(G143), .ZN(new_n901_));
  XNOR2_X1  g765(.A(KEYINPUT54), .B(G132), .ZN(new_n902_));
  AOI22_X1  g766(.A1(new_n628_), .A2(G128), .B1(new_n574_), .B2(new_n902_), .ZN(new_n903_));
  AOI22_X1  g767(.A1(new_n637_), .A2(G159), .B1(new_n552_), .B2(G125), .ZN(new_n904_));
  AOI22_X1  g768(.A1(new_n626_), .A2(G137), .B1(G150), .B2(new_n566_), .ZN(new_n905_));
  AND4_X1   g769(.A1(new_n901_), .A2(new_n903_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g770(.A1(new_n571_), .A2(G124), .ZN(new_n907_));
  XOR2_X1   g771(.A(new_n907_), .B(KEYINPUT55), .Z(new_n908_));
  AOI22_X1  g772(.A1(new_n906_), .A2(new_n908_), .B1(G41), .B2(new_n203_), .ZN(new_n909_));
  AOI21_X1  g773(.A(new_n594_), .B1(new_n900_), .B2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g774(.A(new_n531_), .B1(G50), .B2(new_n825_), .ZN(new_n911_));
  NOR3_X1   g775(.A1(new_n892_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  AND2_X1   g776(.A1(new_n891_), .A2(new_n667_), .ZN(new_n913_));
  AOI22_X1  g777(.A1(new_n654_), .A2(new_n657_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n914_));
  NAND3_X1  g778(.A1(new_n914_), .A2(new_n676_), .A3(new_n606_), .ZN(new_n915_));
  AND3_X1   g779(.A1(new_n914_), .A2(KEYINPUT50), .A3(new_n663_), .ZN(new_n916_));
  AOI21_X1  g780(.A(KEYINPUT50), .B1(new_n914_), .B2(new_n663_), .ZN(new_n917_));
  OAI211_X1 g781(.A(new_n913_), .B(new_n915_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g782(.A(new_n918_), .B1(new_n679_), .B2(new_n891_), .ZN(new_n919_));
  NAND3_X1  g783(.A1(new_n682_), .A2(new_n850_), .A3(G330), .ZN(new_n920_));
  INV_X1    g784(.A(KEYINPUT51), .ZN(new_n921_));
  NAND2_X1  g785(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g786(.A1(new_n525_), .A2(KEYINPUT51), .A3(new_n682_), .ZN(new_n923_));
  AND2_X1   g787(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  OAI21_X1  g788(.A(KEYINPUT52), .B1(new_n919_), .B2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g789(.A1(new_n670_), .A2(KEYINPUT33), .ZN(new_n926_));
  NAND3_X1  g790(.A1(new_n926_), .A2(new_n678_), .A3(new_n658_), .ZN(new_n927_));
  INV_X1    g791(.A(new_n668_), .ZN(new_n928_));
  NAND2_X1  g792(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g793(.A(new_n891_), .ZN(new_n930_));
  NAND2_X1  g794(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g795(.A(KEYINPUT52), .ZN(new_n932_));
  NAND2_X1  g796(.A1(new_n922_), .A2(new_n923_), .ZN(new_n933_));
  NAND4_X1  g797(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .A4(new_n918_), .ZN(new_n934_));
  AOI211_X1 g798(.A(new_n930_), .B(new_n668_), .C1(new_n671_), .C2(new_n678_), .ZN(new_n935_));
  AOI21_X1  g799(.A(new_n891_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n936_));
  OAI21_X1  g800(.A(new_n924_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g801(.A1(new_n925_), .A2(new_n934_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g802(.A(new_n912_), .B1(new_n938_), .B2(new_n530_), .ZN(new_n939_));
  OAI21_X1  g803(.A(new_n865_), .B1(new_n864_), .B2(new_n879_), .ZN(new_n940_));
  NAND3_X1  g804(.A1(new_n931_), .A2(new_n933_), .A3(new_n918_), .ZN(new_n941_));
  NAND2_X1  g805(.A1(new_n919_), .A2(new_n924_), .ZN(new_n942_));
  AOI21_X1  g806(.A(new_n513_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g807(.A1(new_n940_), .A2(new_n943_), .ZN(new_n944_));
  AND2_X1   g808(.A1(new_n939_), .A2(new_n944_), .ZN(new_n945_));
  INV_X1    g809(.A(new_n945_), .ZN(G375));
  OAI211_X1 g810(.A(new_n466_), .B(new_n472_), .C1(new_n526_), .C2(new_n309_), .ZN(new_n947_));
  OAI211_X1 g811(.A(new_n947_), .B(new_n884_), .C1(new_n885_), .C2(new_n844_), .ZN(new_n948_));
  NAND3_X1  g812(.A1(new_n879_), .A2(new_n512_), .A3(new_n948_), .ZN(new_n949_));
  NAND2_X1  g813(.A1(new_n669_), .A2(new_n539_), .ZN(new_n950_));
  OAI21_X1  g814(.A(new_n531_), .B1(G68), .B2(new_n825_), .ZN(new_n951_));
  AOI22_X1  g815(.A1(new_n628_), .A2(G283), .B1(new_n571_), .B2(G303), .ZN(new_n952_));
  OAI21_X1  g816(.A(new_n952_), .B1(new_n335_), .B2(new_n573_), .ZN(new_n953_));
  AOI22_X1  g817(.A1(new_n626_), .A2(G107), .B1(G87), .B2(new_n566_), .ZN(new_n954_));
  AOI22_X1  g818(.A1(G97), .A2(new_n559_), .B1(new_n552_), .B2(G294), .ZN(new_n955_));
  NAND4_X1  g819(.A1(new_n954_), .A2(new_n955_), .A3(G33), .A4(new_n741_), .ZN(new_n956_));
  AOI22_X1  g820(.A1(new_n628_), .A2(G137), .B1(G143), .B2(new_n574_), .ZN(new_n957_));
  NAND2_X1  g821(.A1(new_n571_), .A2(G128), .ZN(new_n958_));
  NAND2_X1  g822(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  AOI22_X1  g823(.A1(new_n626_), .A2(G150), .B1(G50), .B2(new_n566_), .ZN(new_n960_));
  AOI22_X1  g824(.A1(G159), .A2(new_n559_), .B1(new_n552_), .B2(G132), .ZN(new_n961_));
  NAND4_X1  g825(.A1(new_n960_), .A2(new_n961_), .A3(new_n184_), .A4(new_n896_), .ZN(new_n962_));
  OAI22_X1  g826(.A1(new_n953_), .A2(new_n956_), .B1(new_n959_), .B2(new_n962_), .ZN(new_n963_));
  AOI21_X1  g827(.A(new_n951_), .B1(new_n963_), .B2(new_n542_), .ZN(new_n964_));
  AOI22_X1  g828(.A1(new_n886_), .A2(new_n530_), .B1(new_n950_), .B2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g829(.A1(new_n949_), .A2(new_n965_), .ZN(G381));
  INV_X1    g830(.A(G378), .ZN(new_n967_));
  NOR2_X1   g831(.A1(G384), .A2(G381), .ZN(new_n968_));
  NAND3_X1  g832(.A1(new_n945_), .A2(new_n967_), .A3(new_n968_), .ZN(new_n969_));
  OR2_X1    g833(.A1(new_n969_), .A2(KEYINPUT56), .ZN(new_n970_));
  NAND2_X1  g834(.A1(new_n969_), .A2(KEYINPUT56), .ZN(new_n971_));
  NAND4_X1  g835(.A1(new_n733_), .A2(new_n758_), .A3(new_n817_), .A4(new_n823_), .ZN(new_n972_));
  NAND3_X1  g836(.A1(new_n604_), .A2(new_n763_), .A3(new_n789_), .ZN(new_n973_));
  NOR2_X1   g837(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  NAND3_X1  g838(.A1(new_n970_), .A2(new_n971_), .A3(new_n974_), .ZN(new_n975_));
  INV_X1    g839(.A(KEYINPUT57), .ZN(new_n976_));
  XNOR2_X1  g840(.A(new_n975_), .B(new_n976_), .ZN(G407));
  NAND2_X1  g841(.A1(new_n967_), .A2(new_n494_), .ZN(new_n978_));
  INV_X1    g842(.A(new_n978_), .ZN(new_n979_));
  AOI21_X1  g843(.A(new_n491_), .B1(new_n979_), .B2(new_n945_), .ZN(new_n980_));
  NAND2_X1  g844(.A1(G407), .A2(new_n980_), .ZN(G409));
  NAND2_X1  g845(.A1(new_n494_), .A2(G213), .ZN(new_n982_));
  NAND4_X1  g846(.A1(new_n945_), .A2(KEYINPUT58), .A3(G378), .A4(new_n982_), .ZN(new_n983_));
  NAND4_X1  g847(.A1(G378), .A2(new_n939_), .A3(new_n944_), .A4(new_n982_), .ZN(new_n984_));
  INV_X1    g848(.A(KEYINPUT58), .ZN(new_n985_));
  NAND2_X1  g849(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  NAND2_X1  g850(.A1(new_n983_), .A2(new_n986_), .ZN(new_n987_));
  AOI21_X1  g851(.A(new_n865_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n988_));
  NOR2_X1   g852(.A1(new_n864_), .A2(new_n879_), .ZN(new_n989_));
  AOI21_X1  g853(.A(new_n988_), .B1(new_n989_), .B2(new_n938_), .ZN(new_n990_));
  OAI21_X1  g854(.A(new_n939_), .B1(new_n990_), .B2(new_n513_), .ZN(new_n991_));
  OAI211_X1 g855(.A(new_n858_), .B(new_n982_), .C1(new_n880_), .C2(new_n887_), .ZN(new_n992_));
  INV_X1    g856(.A(new_n992_), .ZN(new_n993_));
  NAND2_X1  g857(.A1(new_n991_), .A2(new_n993_), .ZN(new_n994_));
  NAND3_X1  g858(.A1(new_n494_), .A2(G213), .A3(G2897), .ZN(new_n995_));
  INV_X1    g859(.A(new_n995_), .ZN(new_n996_));
  NAND2_X1  g860(.A1(new_n949_), .A2(KEYINPUT59), .ZN(new_n997_));
  INV_X1    g861(.A(KEYINPUT59), .ZN(new_n998_));
  NAND4_X1  g862(.A1(new_n879_), .A2(new_n948_), .A3(new_n998_), .A4(new_n512_), .ZN(new_n999_));
  NAND3_X1  g863(.A1(new_n997_), .A2(new_n965_), .A3(new_n999_), .ZN(new_n1000_));
  AND2_X1   g864(.A1(new_n619_), .A2(new_n645_), .ZN(new_n1001_));
  NAND2_X1  g865(.A1(new_n1000_), .A2(new_n1001_), .ZN(new_n1002_));
  NAND4_X1  g866(.A1(G384), .A2(new_n997_), .A3(new_n965_), .A4(new_n999_), .ZN(new_n1003_));
  AOI21_X1  g867(.A(new_n996_), .B1(new_n1002_), .B2(new_n1003_), .ZN(new_n1004_));
  AND3_X1   g868(.A1(new_n987_), .A2(new_n994_), .A3(new_n1004_), .ZN(new_n1005_));
  NAND2_X1  g869(.A1(new_n1002_), .A2(new_n1003_), .ZN(new_n1006_));
  NAND2_X1  g870(.A1(new_n1006_), .A2(new_n996_), .ZN(new_n1007_));
  AOI21_X1  g871(.A(new_n1007_), .B1(new_n987_), .B2(new_n994_), .ZN(new_n1008_));
  NOR2_X1   g872(.A1(new_n1005_), .A2(new_n1008_), .ZN(new_n1009_));
  NAND2_X1  g873(.A1(G396), .A2(G393), .ZN(new_n1010_));
  AND2_X1   g874(.A1(new_n1010_), .A2(new_n973_), .ZN(new_n1011_));
  AOI21_X1  g875(.A(new_n713_), .B1(new_n529_), .B2(new_n731_), .ZN(new_n1012_));
  INV_X1    g876(.A(new_n758_), .ZN(new_n1013_));
  NOR3_X1   g877(.A1(G390), .A2(new_n1012_), .A3(new_n1013_), .ZN(new_n1014_));
  AOI22_X1  g878(.A1(new_n733_), .A2(new_n758_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n1015_));
  OAI21_X1  g879(.A(new_n1011_), .B1(new_n1014_), .B2(new_n1015_), .ZN(new_n1016_));
  NAND2_X1  g880(.A1(G387), .A2(G390), .ZN(new_n1017_));
  NAND2_X1  g881(.A1(new_n1010_), .A2(new_n973_), .ZN(new_n1018_));
  NAND3_X1  g882(.A1(new_n1017_), .A2(new_n972_), .A3(new_n1018_), .ZN(new_n1019_));
  NAND2_X1  g883(.A1(new_n1016_), .A2(new_n1019_), .ZN(new_n1020_));
  NAND2_X1  g884(.A1(new_n987_), .A2(new_n994_), .ZN(new_n1021_));
  OAI211_X1 g885(.A(new_n1003_), .B(new_n995_), .C1(new_n1002_), .C2(KEYINPUT60), .ZN(new_n1022_));
  AND2_X1   g886(.A1(new_n1002_), .A2(KEYINPUT60), .ZN(new_n1023_));
  NOR2_X1   g887(.A1(new_n1022_), .A2(new_n1023_), .ZN(new_n1024_));
  AOI21_X1  g888(.A(new_n1020_), .B1(new_n1021_), .B2(new_n1024_), .ZN(new_n1025_));
  NAND3_X1  g889(.A1(new_n1002_), .A2(new_n1003_), .A3(new_n996_), .ZN(new_n1026_));
  NAND2_X1  g890(.A1(new_n1026_), .A2(KEYINPUT61), .ZN(new_n1027_));
  INV_X1    g891(.A(KEYINPUT61), .ZN(new_n1028_));
  NAND4_X1  g892(.A1(new_n1002_), .A2(new_n1003_), .A3(new_n1028_), .A4(new_n996_), .ZN(new_n1029_));
  NAND2_X1  g893(.A1(new_n1027_), .A2(new_n1029_), .ZN(new_n1030_));
  AOI22_X1  g894(.A1(new_n983_), .A2(new_n986_), .B1(new_n991_), .B2(new_n993_), .ZN(new_n1031_));
  AOI21_X1  g895(.A(KEYINPUT63), .B1(new_n1030_), .B2(new_n1031_), .ZN(new_n1032_));
  AND3_X1   g896(.A1(new_n1030_), .A2(KEYINPUT63), .A3(new_n1031_), .ZN(new_n1033_));
  OAI211_X1 g897(.A(new_n1009_), .B(new_n1025_), .C1(new_n1032_), .C2(new_n1033_), .ZN(new_n1034_));
  INV_X1    g898(.A(KEYINPUT62), .ZN(new_n1035_));
  NAND3_X1  g899(.A1(new_n1016_), .A2(new_n1019_), .A3(new_n1035_), .ZN(new_n1036_));
  NAND4_X1  g900(.A1(new_n1017_), .A2(new_n1018_), .A3(KEYINPUT62), .A4(new_n972_), .ZN(new_n1037_));
  AND2_X1   g901(.A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1038_));
  NAND2_X1  g902(.A1(new_n1021_), .A2(new_n1024_), .ZN(new_n1039_));
  NAND2_X1  g903(.A1(new_n1030_), .A2(new_n1031_), .ZN(new_n1040_));
  NAND2_X1  g904(.A1(new_n1039_), .A2(new_n1040_), .ZN(new_n1041_));
  NAND3_X1  g905(.A1(new_n987_), .A2(new_n994_), .A3(new_n1004_), .ZN(new_n1042_));
  OAI21_X1  g906(.A(new_n1042_), .B1(new_n1031_), .B2(new_n1007_), .ZN(new_n1043_));
  OAI21_X1  g907(.A(new_n1038_), .B1(new_n1041_), .B2(new_n1043_), .ZN(new_n1044_));
  NAND2_X1  g908(.A1(new_n1034_), .A2(new_n1044_), .ZN(G405));
  XNOR2_X1  g909(.A(new_n945_), .B(G378), .ZN(new_n1046_));
  XNOR2_X1  g910(.A(new_n1046_), .B(new_n1006_), .ZN(new_n1047_));
  NAND2_X1  g911(.A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1048_));
  XNOR2_X1  g912(.A(new_n1047_), .B(new_n1048_), .ZN(G402));
endmodule


