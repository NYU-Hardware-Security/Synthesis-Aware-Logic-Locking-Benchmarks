//Secret key is'1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_c6288" written by ABC on Sun Nov 20 19:50:26 2022

module locked_c6288 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1gat, G18gat, G35gat, G52gat, G69gat,
    G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat,
    G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat,
    G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat,
    G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1gat, G18gat, G35gat, G52gat,
    G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat,
    G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat,
    G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat,
    G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_n193_, new_n194_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_,
    new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_,
    new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_,
    new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_,
    new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_,
    new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2949_, new_n2950_;
  INV_X1    g0000(.A(G1gat), .ZN(new_n193_));
  INV_X1    g0001(.A(G273gat), .ZN(new_n194_));
  NOR2_X1   g0002(.A1(new_n193_), .A2(new_n194_), .ZN(G545gat));
  INV_X1    g0003(.A(G18gat), .ZN(new_n196_));
  NOR2_X1   g0004(.A1(new_n196_), .A2(new_n194_), .ZN(new_n197_));
  INV_X1    g0005(.A(G290gat), .ZN(new_n198_));
  NOR2_X1   g0006(.A1(new_n193_), .A2(new_n198_), .ZN(new_n199_));
  NAND2_X1  g0007(.A1(new_n197_), .A2(new_n199_), .ZN(new_n200_));
  INV_X1    g0008(.A(new_n200_), .ZN(new_n201_));
  NOR2_X1   g0009(.A1(new_n197_), .A2(new_n199_), .ZN(new_n202_));
  NOR2_X1   g0010(.A1(new_n201_), .A2(new_n202_), .ZN(G1581gat));
  NAND3_X1  g0011(.A1(new_n197_), .A2(G35gat), .A3(G290gat), .ZN(new_n204_));
  INV_X1    g0012(.A(G35gat), .ZN(new_n205_));
  OAI22_X1  g0013(.A1(new_n196_), .A2(new_n198_), .B1(new_n205_), .B2(new_n194_), .ZN(new_n206_));
  NAND3_X1  g0014(.A1(new_n204_), .A2(KEYINPUT0), .A3(new_n206_), .ZN(new_n207_));
  OAI211_X1 g0015(.A(new_n207_), .B(new_n200_), .C1(KEYINPUT0), .C2(new_n206_), .ZN(new_n208_));
  NAND3_X1  g0016(.A1(new_n201_), .A2(KEYINPUT0), .A3(new_n204_), .ZN(new_n209_));
  NAND2_X1  g0017(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g0018(.A(G307gat), .ZN(new_n211_));
  NOR2_X1   g0019(.A1(new_n193_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g0020(.A(new_n210_), .B(new_n212_), .ZN(G1901gat));
  INV_X1    g0021(.A(new_n204_), .ZN(new_n214_));
  INV_X1    g0022(.A(G52gat), .ZN(new_n215_));
  OAI22_X1  g0023(.A1(new_n205_), .A2(new_n198_), .B1(new_n215_), .B2(new_n194_), .ZN(new_n216_));
  NAND4_X1  g0024(.A1(G35gat), .A2(G52gat), .A3(G273gat), .A4(G290gat), .ZN(new_n217_));
  NAND2_X1  g0025(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g0026(.A1(new_n218_), .A2(KEYINPUT1), .ZN(new_n219_));
  INV_X1    g0027(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g0028(.A1(new_n218_), .A2(KEYINPUT1), .ZN(new_n221_));
  AOI21_X1  g0029(.A(new_n214_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g0030(.A1(new_n219_), .A2(new_n204_), .ZN(new_n223_));
  OR4_X1    g0031(.A1(new_n196_), .A2(new_n222_), .A3(new_n211_), .A4(new_n223_), .ZN(new_n224_));
  OAI22_X1  g0032(.A1(new_n222_), .A2(new_n223_), .B1(new_n196_), .B2(new_n211_), .ZN(new_n225_));
  AND2_X1   g0033(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g0034(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n227_));
  NAND2_X1  g0035(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g0036(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g0037(.A1(new_n226_), .A2(new_n227_), .ZN(new_n230_));
  NOR2_X1   g0038(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g0039(.A(G324gat), .ZN(new_n232_));
  NOR2_X1   g0040(.A1(new_n193_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g0041(.A(new_n231_), .B(new_n233_), .Z(G2223gat));
  NAND2_X1  g0042(.A1(new_n218_), .A2(new_n204_), .ZN(new_n235_));
  XNOR2_X1  g0043(.A(new_n235_), .B(KEYINPUT2), .ZN(new_n236_));
  NAND2_X1  g0044(.A1(new_n225_), .A2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g0045(.A1(G52gat), .A2(G69gat), .A3(G273gat), .A4(G290gat), .ZN(new_n238_));
  INV_X1    g0046(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g0047(.A1(new_n239_), .A2(new_n217_), .ZN(new_n240_));
  INV_X1    g0048(.A(G69gat), .ZN(new_n241_));
  OAI22_X1  g0049(.A1(new_n215_), .A2(new_n198_), .B1(new_n241_), .B2(new_n194_), .ZN(new_n242_));
  NAND2_X1  g0050(.A1(new_n242_), .A2(new_n238_), .ZN(new_n243_));
  AOI21_X1  g0051(.A(new_n240_), .B1(new_n217_), .B2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g0052(.A1(new_n205_), .A2(new_n211_), .ZN(new_n245_));
  XNOR2_X1  g0053(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g0054(.A1(new_n237_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g0055(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g0056(.A1(new_n237_), .A2(new_n246_), .ZN(new_n249_));
  NOR2_X1   g0057(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g0058(.A1(new_n196_), .A2(new_n232_), .ZN(new_n251_));
  XNOR2_X1  g0059(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  OAI21_X1  g0060(.A(new_n228_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n253_));
  NAND2_X1  g0061(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g0062(.A(new_n254_), .ZN(new_n255_));
  NOR2_X1   g0063(.A1(new_n252_), .A2(new_n253_), .ZN(new_n256_));
  NOR2_X1   g0064(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g0065(.A(G341gat), .ZN(new_n258_));
  NOR2_X1   g0066(.A1(new_n193_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g0067(.A(new_n257_), .B(new_n259_), .Z(G2548gat));
  OAI21_X1  g0068(.A(new_n254_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n261_));
  OAI21_X1  g0069(.A(new_n247_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n262_));
  NAND4_X1  g0070(.A1(G69gat), .A2(G86gat), .A3(G273gat), .A4(G290gat), .ZN(new_n263_));
  INV_X1    g0071(.A(new_n263_), .ZN(new_n264_));
  AOI22_X1  g0072(.A1(G69gat), .A2(G290gat), .B1(G86gat), .B2(G273gat), .ZN(new_n265_));
  OAI21_X1  g0073(.A(new_n238_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g0074(.A1(new_n239_), .A2(new_n263_), .ZN(new_n267_));
  NAND2_X1  g0075(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g0076(.A1(G52gat), .A2(G307gat), .ZN(new_n269_));
  XNOR2_X1  g0077(.A(new_n269_), .B(KEYINPUT3), .ZN(new_n270_));
  XNOR2_X1  g0078(.A(new_n268_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g0079(.A1(new_n243_), .A2(new_n217_), .ZN(new_n272_));
  OAI21_X1  g0080(.A(new_n272_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n273_));
  NOR2_X1   g0081(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g0082(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g0083(.A1(new_n271_), .A2(new_n273_), .ZN(new_n276_));
  NAND2_X1  g0084(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g0085(.A1(new_n205_), .A2(new_n232_), .ZN(new_n278_));
  INV_X1    g0086(.A(KEYINPUT4), .ZN(new_n279_));
  XNOR2_X1  g0087(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g0088(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g0089(.A(new_n275_), .B(new_n276_), .C1(new_n279_), .C2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g0090(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g0091(.A1(new_n262_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g0092(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g0093(.A1(G18gat), .A2(G341gat), .ZN(new_n286_));
  NAND2_X1  g0094(.A1(new_n262_), .A2(new_n283_), .ZN(new_n287_));
  NAND3_X1  g0095(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g0096(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g0097(.A(new_n286_), .B1(new_n287_), .B2(new_n285_), .ZN(new_n290_));
  NOR2_X1   g0098(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g0099(.A1(new_n261_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g0100(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g0101(.A1(new_n261_), .A2(new_n291_), .ZN(new_n294_));
  NOR2_X1   g0102(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g0103(.A1(KEYINPUT5), .A2(G358gat), .ZN(new_n296_));
  INV_X1    g0104(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g0105(.A1(KEYINPUT5), .A2(G358gat), .ZN(new_n298_));
  NOR2_X1   g0106(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g0107(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g0108(.A1(new_n300_), .A2(new_n193_), .ZN(new_n301_));
  INV_X1    g0109(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g0110(.A(new_n295_), .B(new_n302_), .ZN(G2877gat));
  OAI21_X1  g0111(.A(new_n292_), .B1(new_n294_), .B2(new_n301_), .ZN(new_n304_));
  NOR2_X1   g0112(.A1(new_n215_), .A2(new_n232_), .ZN(new_n305_));
  INV_X1    g0113(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g0114(.A1(new_n266_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n307_));
  NAND2_X1  g0115(.A1(new_n307_), .A2(new_n266_), .ZN(new_n308_));
  NAND2_X1  g0116(.A1(G103gat), .A2(G290gat), .ZN(new_n309_));
  INV_X1    g0117(.A(G86gat), .ZN(new_n310_));
  NOR3_X1   g0118(.A1(new_n309_), .A2(new_n310_), .A3(new_n194_), .ZN(new_n311_));
  NOR2_X1   g0119(.A1(new_n311_), .A2(new_n263_), .ZN(new_n312_));
  INV_X1    g0120(.A(new_n312_), .ZN(new_n313_));
  AND2_X1   g0121(.A1(G103gat), .A2(G290gat), .ZN(new_n314_));
  NAND3_X1  g0122(.A1(new_n314_), .A2(G86gat), .A3(G273gat), .ZN(new_n315_));
  NAND2_X1  g0123(.A1(G103gat), .A2(G273gat), .ZN(new_n316_));
  OAI21_X1  g0124(.A(new_n316_), .B1(new_n310_), .B2(new_n198_), .ZN(new_n317_));
  NAND2_X1  g0125(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g0126(.A1(new_n318_), .A2(new_n263_), .ZN(new_n319_));
  NAND2_X1  g0127(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g0128(.A1(G69gat), .A2(G307gat), .ZN(new_n321_));
  INV_X1    g0129(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g0130(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g0131(.A1(new_n313_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n324_));
  AOI21_X1  g0132(.A(new_n308_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g0133(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g0134(.A1(new_n323_), .A2(new_n308_), .A3(new_n324_), .ZN(new_n327_));
  AOI21_X1  g0135(.A(new_n306_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g0136(.A1(new_n276_), .A2(new_n278_), .ZN(new_n329_));
  NAND2_X1  g0137(.A1(new_n329_), .A2(new_n275_), .ZN(new_n330_));
  INV_X1    g0138(.A(new_n327_), .ZN(new_n331_));
  NOR3_X1   g0139(.A1(new_n331_), .A2(new_n325_), .A3(new_n305_), .ZN(new_n332_));
  NOR3_X1   g0140(.A1(new_n328_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g0141(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g0142(.A1(new_n205_), .A2(new_n258_), .ZN(new_n335_));
  INV_X1    g0143(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g0144(.A(new_n330_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n337_));
  NAND3_X1  g0145(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g0146(.A(new_n337_), .ZN(new_n339_));
  OAI21_X1  g0147(.A(new_n335_), .B1(new_n339_), .B2(new_n333_), .ZN(new_n340_));
  AND2_X1   g0148(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g0149(.A1(new_n288_), .A2(KEYINPUT6), .ZN(new_n342_));
  INV_X1    g0150(.A(new_n287_), .ZN(new_n343_));
  AOI21_X1  g0151(.A(new_n343_), .B1(new_n288_), .B2(KEYINPUT6), .ZN(new_n344_));
  AOI21_X1  g0152(.A(new_n341_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g0153(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g0154(.A1(new_n341_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n347_));
  NAND4_X1  g0155(.A1(new_n346_), .A2(G18gat), .A3(new_n299_), .A4(new_n347_), .ZN(new_n348_));
  INV_X1    g0156(.A(new_n347_), .ZN(new_n349_));
  OAI22_X1  g0157(.A1(new_n345_), .A2(new_n349_), .B1(new_n196_), .B2(new_n300_), .ZN(new_n350_));
  AOI21_X1  g0158(.A(new_n304_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g0159(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g0160(.A1(new_n348_), .A2(new_n304_), .A3(new_n350_), .ZN(new_n353_));
  NAND2_X1  g0161(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g0162(.A(G375gat), .ZN(new_n355_));
  NOR2_X1   g0163(.A1(new_n193_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g0164(.A(new_n354_), .B(new_n356_), .ZN(G3211gat));
  NOR2_X1   g0165(.A1(new_n196_), .A2(new_n355_), .ZN(new_n358_));
  NAND2_X1  g0166(.A1(new_n342_), .A2(new_n344_), .ZN(new_n359_));
  NAND2_X1  g0167(.A1(new_n359_), .A2(new_n341_), .ZN(new_n360_));
  NOR2_X1   g0168(.A1(new_n300_), .A2(new_n205_), .ZN(new_n361_));
  AOI21_X1  g0169(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n362_));
  NAND2_X1  g0170(.A1(G69gat), .A2(G324gat), .ZN(new_n363_));
  NAND4_X1  g0171(.A1(G103gat), .A2(G120gat), .A3(G273gat), .A4(G290gat), .ZN(new_n364_));
  INV_X1    g0172(.A(new_n364_), .ZN(new_n365_));
  AOI22_X1  g0173(.A1(G103gat), .A2(G290gat), .B1(G120gat), .B2(G273gat), .ZN(new_n366_));
  OAI21_X1  g0174(.A(new_n315_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g0175(.A1(new_n364_), .A2(new_n314_), .A3(G86gat), .A4(G273gat), .ZN(new_n368_));
  NAND2_X1  g0176(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g0177(.A1(G86gat), .A2(G307gat), .ZN(new_n370_));
  NAND3_X1  g0178(.A1(new_n369_), .A2(KEYINPUT7), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g0179(.A(new_n319_), .B1(new_n312_), .B2(new_n322_), .ZN(new_n372_));
  NAND2_X1  g0180(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g0181(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n375_));
  INV_X1    g0183(.A(new_n316_), .ZN(new_n376_));
  AND2_X1   g0184(.A1(G120gat), .A2(G290gat), .ZN(new_n377_));
  NAND2_X1  g0185(.A1(G120gat), .A2(G273gat), .ZN(new_n378_));
  AOI22_X1  g0186(.A1(new_n376_), .A2(new_n377_), .B1(new_n309_), .B2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g0187(.A(new_n370_), .B(new_n368_), .C1(new_n379_), .C2(new_n311_), .ZN(new_n380_));
  INV_X1    g0188(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g0189(.A(new_n370_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n382_));
  OAI21_X1  g0190(.A(new_n375_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g0191(.A1(new_n374_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g0192(.A(new_n324_), .B(new_n319_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n385_));
  AOI21_X1  g0193(.A(new_n363_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g0194(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g0195(.A(new_n327_), .B1(new_n325_), .B2(new_n305_), .ZN(new_n388_));
  INV_X1    g0196(.A(new_n383_), .ZN(new_n389_));
  OAI211_X1 g0197(.A(new_n385_), .B(new_n363_), .C1(new_n389_), .C2(new_n373_), .ZN(new_n390_));
  NAND3_X1  g0198(.A1(new_n387_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  NOR2_X1   g0199(.A1(new_n215_), .A2(new_n258_), .ZN(new_n392_));
  INV_X1    g0200(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g0201(.A(new_n388_), .ZN(new_n394_));
  INV_X1    g0202(.A(new_n390_), .ZN(new_n395_));
  OAI21_X1  g0203(.A(new_n394_), .B1(new_n395_), .B2(new_n386_), .ZN(new_n396_));
  NAND3_X1  g0204(.A1(new_n391_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g0205(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g0206(.A(new_n393_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g0207(.A(new_n362_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g0208(.A(new_n400_), .ZN(new_n401_));
  NOR3_X1   g0209(.A1(new_n398_), .A2(new_n362_), .A3(new_n399_), .ZN(new_n402_));
  OAI21_X1  g0210(.A(new_n361_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g0211(.A(new_n362_), .ZN(new_n404_));
  INV_X1    g0212(.A(new_n399_), .ZN(new_n405_));
  NAND3_X1  g0213(.A1(new_n404_), .A2(new_n397_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g0214(.A(new_n361_), .ZN(new_n407_));
  NAND3_X1  g0215(.A1(new_n406_), .A2(new_n407_), .A3(new_n400_), .ZN(new_n408_));
  NAND2_X1  g0216(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  AND3_X1   g0217(.A1(new_n350_), .A2(new_n360_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g0218(.A(new_n409_), .B1(new_n350_), .B2(new_n360_), .ZN(new_n411_));
  OAI21_X1  g0219(.A(new_n358_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g0220(.A1(new_n350_), .A2(new_n360_), .ZN(new_n413_));
  INV_X1    g0221(.A(new_n409_), .ZN(new_n414_));
  NAND2_X1  g0222(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g0223(.A(new_n358_), .ZN(new_n416_));
  NAND3_X1  g0224(.A1(new_n350_), .A2(new_n360_), .A3(new_n409_), .ZN(new_n417_));
  NAND3_X1  g0225(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g0226(.A1(new_n412_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g0227(.A(new_n353_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n420_));
  INV_X1    g0228(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g0229(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g0230(.A1(new_n420_), .A2(new_n418_), .A3(new_n412_), .ZN(new_n423_));
  NAND2_X1  g0231(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g0232(.A1(G1gat), .A2(G392gat), .ZN(new_n425_));
  XOR2_X1   g0233(.A(new_n425_), .B(KEYINPUT8), .Z(new_n426_));
  XOR2_X1   g0234(.A(new_n424_), .B(new_n426_), .Z(G3552gat));
  INV_X1    g0235(.A(new_n423_), .ZN(new_n428_));
  OR2_X1    g0236(.A1(new_n428_), .A2(KEYINPUT9), .ZN(new_n429_));
  NAND3_X1  g0237(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n430_));
  NAND2_X1  g0238(.A1(new_n428_), .A2(KEYINPUT9), .ZN(new_n431_));
  NAND3_X1  g0239(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g0240(.A(new_n411_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n433_));
  AOI21_X1  g0241(.A(new_n402_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n434_));
  INV_X1    g0242(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g0243(.A1(new_n300_), .A2(new_n215_), .ZN(new_n436_));
  INV_X1    g0244(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g0245(.A(KEYINPUT11), .ZN(new_n438_));
  NAND2_X1  g0246(.A1(new_n397_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g0247(.A1(new_n310_), .A2(new_n232_), .ZN(new_n440_));
  INV_X1    g0248(.A(KEYINPUT12), .ZN(new_n441_));
  OAI21_X1  g0249(.A(new_n441_), .B1(new_n379_), .B2(new_n311_), .ZN(new_n442_));
  OAI211_X1 g0250(.A(new_n315_), .B(KEYINPUT12), .C1(new_n365_), .C2(new_n366_), .ZN(new_n443_));
  AND3_X1   g0251(.A1(new_n380_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g0252(.A1(G120gat), .A2(G290gat), .ZN(new_n445_));
  NAND2_X1  g0253(.A1(G137gat), .A2(G273gat), .ZN(new_n446_));
  NAND2_X1  g0254(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g0255(.A1(G120gat), .A2(G137gat), .A3(G273gat), .A4(G290gat), .ZN(new_n448_));
  AOI22_X1  g0256(.A1(new_n447_), .A2(new_n448_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n449_));
  AND4_X1   g0257(.A1(G120gat), .A2(G137gat), .A3(G273gat), .A4(G290gat), .ZN(new_n450_));
  NOR2_X1   g0258(.A1(new_n450_), .A2(new_n364_), .ZN(new_n451_));
  INV_X1    g0259(.A(G103gat), .ZN(new_n452_));
  NOR2_X1   g0260(.A1(new_n452_), .A2(new_n211_), .ZN(new_n453_));
  NOR3_X1   g0261(.A1(new_n449_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g0262(.A(new_n453_), .ZN(new_n455_));
  AOI22_X1  g0263(.A1(G120gat), .A2(G290gat), .B1(G137gat), .B2(G273gat), .ZN(new_n456_));
  OAI21_X1  g0264(.A(new_n364_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g0265(.A1(new_n365_), .A2(new_n448_), .ZN(new_n458_));
  AOI21_X1  g0266(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g0267(.A(KEYINPUT13), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g0268(.A(new_n453_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n461_));
  NAND3_X1  g0269(.A1(new_n457_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n462_));
  INV_X1    g0270(.A(KEYINPUT13), .ZN(new_n463_));
  NAND3_X1  g0271(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g0272(.A(new_n444_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g0273(.A(new_n463_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n466_));
  NAND3_X1  g0274(.A1(new_n380_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n467_));
  NOR2_X1   g0275(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g0276(.A(new_n440_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g0277(.A(KEYINPUT14), .ZN(new_n470_));
  AND3_X1   g0278(.A1(new_n461_), .A2(new_n463_), .A3(new_n462_), .ZN(new_n471_));
  OAI21_X1  g0279(.A(new_n467_), .B1(new_n471_), .B2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g0280(.A1(new_n460_), .A2(new_n444_), .ZN(new_n473_));
  INV_X1    g0281(.A(new_n440_), .ZN(new_n474_));
  NAND3_X1  g0282(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g0283(.A1(new_n469_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  NAND4_X1  g0284(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT14), .A4(new_n474_), .ZN(new_n477_));
  NAND2_X1  g0285(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI22_X1  g0286(.A1(new_n374_), .A2(new_n383_), .B1(new_n385_), .B2(new_n363_), .ZN(new_n479_));
  NAND2_X1  g0287(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g0288(.A1(new_n241_), .A2(new_n258_), .ZN(new_n481_));
  INV_X1    g0289(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g0290(.A(new_n479_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n483_));
  INV_X1    g0291(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g0292(.A1(new_n480_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g0293(.A(new_n479_), .ZN(new_n486_));
  AOI21_X1  g0294(.A(new_n486_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n487_));
  OAI21_X1  g0295(.A(new_n481_), .B1(new_n487_), .B2(new_n483_), .ZN(new_n488_));
  NAND3_X1  g0296(.A1(new_n439_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g0297(.A(KEYINPUT10), .ZN(new_n490_));
  NAND2_X1  g0298(.A1(new_n391_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g0299(.A1(new_n387_), .A2(new_n388_), .A3(KEYINPUT10), .A4(new_n390_), .ZN(new_n492_));
  NAND3_X1  g0300(.A1(new_n397_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g0301(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g0302(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g0303(.A1(new_n493_), .A2(new_n439_), .A3(new_n485_), .A4(new_n488_), .ZN(new_n496_));
  AOI21_X1  g0304(.A(new_n437_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g0305(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g0306(.A1(new_n495_), .A2(new_n437_), .A3(new_n496_), .ZN(new_n499_));
  AOI21_X1  g0307(.A(new_n435_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g0308(.A(new_n499_), .ZN(new_n501_));
  NOR3_X1   g0309(.A1(new_n501_), .A2(new_n434_), .A3(new_n497_), .ZN(new_n502_));
  NOR2_X1   g0310(.A1(new_n205_), .A2(new_n355_), .ZN(new_n503_));
  NOR3_X1   g0311(.A1(new_n500_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g0312(.A(new_n503_), .ZN(new_n505_));
  OAI21_X1  g0313(.A(new_n434_), .B1(new_n501_), .B2(new_n497_), .ZN(new_n506_));
  NAND3_X1  g0314(.A1(new_n498_), .A2(new_n435_), .A3(new_n499_), .ZN(new_n507_));
  AOI21_X1  g0315(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g0316(.A(new_n433_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g0317(.A(new_n415_), .B1(new_n410_), .B2(new_n358_), .ZN(new_n510_));
  NOR2_X1   g0318(.A1(new_n504_), .A2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g0319(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g0320(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g0321(.A1(G18gat), .A2(G392gat), .ZN(new_n514_));
  XNOR2_X1  g0322(.A(new_n514_), .B(KEYINPUT15), .ZN(new_n515_));
  NAND2_X1  g0323(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g0324(.A(new_n515_), .ZN(new_n517_));
  NAND3_X1  g0325(.A1(new_n509_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g0326(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g0327(.A1(new_n432_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g0328(.A1(new_n422_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n521_));
  NAND3_X1  g0329(.A1(new_n429_), .A2(new_n521_), .A3(new_n431_), .ZN(new_n522_));
  OAI21_X1  g0330(.A(new_n520_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g0331(.A1(G1gat), .A2(G409gat), .ZN(new_n524_));
  XNOR2_X1  g0332(.A(new_n523_), .B(new_n524_), .ZN(G3895gat));
  NAND2_X1  g0333(.A1(new_n523_), .A2(new_n524_), .ZN(new_n526_));
  NAND3_X1  g0334(.A1(new_n432_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n527_));
  NAND2_X1  g0335(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g0336(.A(new_n507_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n529_));
  NOR2_X1   g0337(.A1(new_n452_), .A2(new_n232_), .ZN(new_n530_));
  INV_X1    g0338(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g0339(.A(G120gat), .ZN(new_n532_));
  NOR2_X1   g0340(.A1(new_n532_), .A2(new_n211_), .ZN(new_n533_));
  NAND2_X1  g0341(.A1(G137gat), .A2(G290gat), .ZN(new_n534_));
  NAND2_X1  g0342(.A1(G154gat), .A2(G273gat), .ZN(new_n535_));
  NAND2_X1  g0343(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g0344(.A1(G137gat), .A2(G154gat), .A3(G273gat), .A4(G290gat), .ZN(new_n537_));
  INV_X1    g0345(.A(new_n378_), .ZN(new_n538_));
  AND2_X1   g0346(.A1(G137gat), .A2(G290gat), .ZN(new_n539_));
  AOI22_X1  g0347(.A1(new_n536_), .A2(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND4_X1   g0348(.A1(G137gat), .A2(G154gat), .A3(G273gat), .A4(G290gat), .ZN(new_n541_));
  NOR2_X1   g0349(.A1(new_n541_), .A2(new_n448_), .ZN(new_n542_));
  OAI21_X1  g0350(.A(new_n533_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  AOI22_X1  g0351(.A1(G137gat), .A2(G290gat), .B1(G154gat), .B2(G273gat), .ZN(new_n544_));
  OAI21_X1  g0352(.A(new_n448_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g0353(.A(new_n533_), .ZN(new_n546_));
  NAND2_X1  g0354(.A1(new_n450_), .A2(new_n537_), .ZN(new_n547_));
  NAND3_X1  g0355(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g0356(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g0357(.A(KEYINPUT17), .ZN(new_n550_));
  OAI211_X1 g0358(.A(new_n457_), .B(new_n550_), .C1(new_n453_), .C2(new_n451_), .ZN(new_n551_));
  OAI21_X1  g0359(.A(new_n457_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n552_));
  NAND2_X1  g0360(.A1(new_n552_), .A2(KEYINPUT17), .ZN(new_n553_));
  AOI21_X1  g0361(.A(new_n549_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  AND2_X1   g0362(.A1(new_n549_), .A2(new_n551_), .ZN(new_n555_));
  OAI21_X1  g0363(.A(new_n531_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g0364(.A1(new_n553_), .A2(new_n551_), .ZN(new_n557_));
  INV_X1    g0365(.A(new_n549_), .ZN(new_n558_));
  NAND2_X1  g0366(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g0367(.A1(new_n549_), .A2(new_n551_), .ZN(new_n560_));
  NAND3_X1  g0368(.A1(new_n559_), .A2(new_n530_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g0369(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g0370(.A(new_n474_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n563_));
  NOR3_X1   g0371(.A1(new_n444_), .A2(new_n454_), .A3(new_n459_), .ZN(new_n564_));
  INV_X1    g0372(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g0373(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g0374(.A(new_n440_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n567_));
  OAI211_X1 g0375(.A(new_n556_), .B(new_n561_), .C1(new_n567_), .C2(new_n564_), .ZN(new_n568_));
  NAND2_X1  g0376(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g0377(.A1(new_n310_), .A2(new_n258_), .ZN(new_n570_));
  NAND2_X1  g0378(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g0379(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g0380(.A1(new_n566_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g0381(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g0382(.A1(new_n487_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n575_));
  NOR2_X1   g0383(.A1(new_n478_), .A2(new_n479_), .ZN(new_n576_));
  OAI21_X1  g0384(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g0385(.A(new_n576_), .ZN(new_n578_));
  NAND4_X1  g0386(.A1(new_n485_), .A2(new_n578_), .A3(new_n573_), .A4(new_n571_), .ZN(new_n579_));
  NAND2_X1  g0387(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g0388(.A1(new_n300_), .A2(new_n241_), .ZN(new_n581_));
  INV_X1    g0389(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g0390(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g0391(.A(new_n581_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n584_));
  NOR2_X1   g0392(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g0393(.A1(new_n493_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n586_));
  NAND2_X1  g0394(.A1(new_n499_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g0395(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g0396(.A1(new_n215_), .A2(new_n355_), .ZN(new_n589_));
  INV_X1    g0397(.A(new_n589_), .ZN(new_n590_));
  OAI211_X1 g0398(.A(new_n499_), .B(new_n586_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n591_));
  NAND3_X1  g0399(.A1(new_n588_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g0400(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g0401(.A(new_n590_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n594_));
  OAI21_X1  g0402(.A(new_n529_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g0403(.A1(new_n588_), .A2(new_n591_), .ZN(new_n596_));
  NAND2_X1  g0404(.A1(new_n596_), .A2(new_n589_), .ZN(new_n597_));
  AOI21_X1  g0405(.A(new_n502_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n598_));
  NAND3_X1  g0406(.A1(new_n597_), .A2(new_n598_), .A3(new_n592_), .ZN(new_n599_));
  NAND2_X1  g0407(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g0408(.A(G392gat), .ZN(new_n601_));
  NOR2_X1   g0409(.A1(new_n205_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g0410(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g0411(.A(new_n600_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g0412(.A(KEYINPUT18), .ZN(new_n605_));
  NAND2_X1  g0413(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g0414(.A1(new_n513_), .A2(KEYINPUT16), .ZN(new_n607_));
  INV_X1    g0415(.A(KEYINPUT16), .ZN(new_n608_));
  NAND3_X1  g0416(.A1(new_n509_), .A2(new_n512_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g0417(.A1(new_n607_), .A2(new_n517_), .A3(new_n609_), .ZN(new_n610_));
  NAND4_X1  g0418(.A1(new_n595_), .A2(new_n599_), .A3(KEYINPUT18), .A4(new_n603_), .ZN(new_n611_));
  NAND4_X1  g0419(.A1(new_n606_), .A2(new_n610_), .A3(new_n512_), .A4(new_n611_), .ZN(new_n612_));
  INV_X1    g0420(.A(G409gat), .ZN(new_n613_));
  NOR2_X1   g0421(.A1(new_n196_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g0422(.A1(new_n512_), .A2(G18gat), .A3(G392gat), .ZN(new_n615_));
  AND2_X1   g0423(.A1(new_n615_), .A2(new_n509_), .ZN(new_n616_));
  NAND2_X1  g0424(.A1(new_n616_), .A2(new_n604_), .ZN(new_n617_));
  AND3_X1   g0425(.A1(new_n612_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g0426(.A(new_n614_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g0427(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OR2_X1    g0428(.A1(new_n528_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g0429(.A1(new_n528_), .A2(new_n620_), .ZN(new_n622_));
  NAND2_X1  g0430(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g0431(.A(G426gat), .ZN(new_n624_));
  NOR2_X1   g0432(.A1(new_n193_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g0433(.A(new_n623_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g0434(.A(new_n626_), .B(KEYINPUT19), .ZN(G4241gat));
  INV_X1    g0435(.A(new_n622_), .ZN(new_n628_));
  INV_X1    g0436(.A(new_n625_), .ZN(new_n629_));
  AOI21_X1  g0437(.A(new_n628_), .B1(new_n621_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g0438(.A(new_n619_), .ZN(new_n631_));
  AND2_X1   g0439(.A1(new_n606_), .A2(new_n611_), .ZN(new_n632_));
  NAND2_X1  g0440(.A1(new_n632_), .A2(new_n616_), .ZN(new_n633_));
  NOR2_X1   g0441(.A1(new_n205_), .A2(new_n613_), .ZN(new_n634_));
  INV_X1    g0442(.A(KEYINPUT20), .ZN(new_n635_));
  OAI21_X1  g0443(.A(new_n635_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n636_));
  NAND3_X1  g0444(.A1(new_n597_), .A2(KEYINPUT20), .A3(new_n592_), .ZN(new_n637_));
  NAND3_X1  g0445(.A1(new_n636_), .A2(new_n637_), .A3(new_n529_), .ZN(new_n638_));
  AOI21_X1  g0446(.A(new_n602_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n639_));
  OAI21_X1  g0447(.A(new_n638_), .B1(new_n639_), .B2(KEYINPUT29), .ZN(new_n640_));
  AND3_X1   g0448(.A1(new_n600_), .A2(KEYINPUT29), .A3(new_n603_), .ZN(new_n641_));
  NAND2_X1  g0449(.A1(G69gat), .A2(G375gat), .ZN(new_n642_));
  XOR2_X1   g0450(.A(new_n642_), .B(KEYINPUT28), .Z(new_n643_));
  INV_X1    g0451(.A(new_n568_), .ZN(new_n644_));
  AOI21_X1  g0452(.A(new_n644_), .B1(new_n572_), .B2(new_n566_), .ZN(new_n645_));
  NAND2_X1  g0453(.A1(new_n558_), .A2(new_n552_), .ZN(new_n646_));
  AND2_X1   g0454(.A1(new_n556_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g0455(.A1(new_n532_), .A2(new_n232_), .ZN(new_n648_));
  INV_X1    g0456(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g0457(.A(KEYINPUT25), .ZN(new_n650_));
  INV_X1    g0458(.A(G137gat), .ZN(new_n651_));
  NOR2_X1   g0459(.A1(new_n651_), .A2(new_n211_), .ZN(new_n652_));
  INV_X1    g0460(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g0461(.A1(G154gat), .A2(G290gat), .ZN(new_n654_));
  NAND2_X1  g0462(.A1(G171gat), .A2(G273gat), .ZN(new_n655_));
  NAND2_X1  g0463(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g0464(.A1(G154gat), .A2(G171gat), .A3(G273gat), .A4(G290gat), .ZN(new_n657_));
  AND2_X1   g0465(.A1(G137gat), .A2(G273gat), .ZN(new_n658_));
  AND2_X1   g0466(.A1(G154gat), .A2(G290gat), .ZN(new_n659_));
  AOI22_X1  g0467(.A1(new_n656_), .A2(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AND4_X1   g0468(.A1(G154gat), .A2(G171gat), .A3(G273gat), .A4(G290gat), .ZN(new_n661_));
  NOR2_X1   g0469(.A1(new_n661_), .A2(new_n537_), .ZN(new_n662_));
  OAI21_X1  g0470(.A(new_n653_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  AOI22_X1  g0471(.A1(G154gat), .A2(G290gat), .B1(G171gat), .B2(G273gat), .ZN(new_n664_));
  OAI21_X1  g0472(.A(new_n537_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g0473(.A1(new_n541_), .A2(new_n657_), .ZN(new_n666_));
  NAND3_X1  g0474(.A1(new_n665_), .A2(new_n652_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g0475(.A(new_n650_), .B1(new_n663_), .B2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g0476(.A1(new_n660_), .A2(new_n662_), .ZN(new_n669_));
  AOI21_X1  g0477(.A(KEYINPUT25), .B1(new_n669_), .B2(new_n652_), .ZN(new_n670_));
  AOI21_X1  g0478(.A(new_n540_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n671_));
  NOR3_X1   g0479(.A1(new_n668_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n673_));
  NAND2_X1  g0481(.A1(new_n545_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g0482(.A1(new_n540_), .A2(KEYINPUT26), .ZN(new_n675_));
  NAND3_X1  g0483(.A1(new_n548_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g0484(.A(new_n676_), .B1(new_n663_), .B2(new_n667_), .ZN(new_n677_));
  OAI21_X1  g0485(.A(new_n649_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g0486(.A1(new_n663_), .A2(new_n667_), .ZN(new_n679_));
  NAND2_X1  g0487(.A1(new_n679_), .A2(KEYINPUT25), .ZN(new_n680_));
  INV_X1    g0488(.A(new_n671_), .ZN(new_n681_));
  NAND2_X1  g0489(.A1(new_n667_), .A2(new_n650_), .ZN(new_n682_));
  NAND3_X1  g0490(.A1(new_n680_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  NAND4_X1  g0491(.A1(new_n679_), .A2(new_n548_), .A3(new_n674_), .A4(new_n675_), .ZN(new_n684_));
  NAND3_X1  g0492(.A1(new_n683_), .A2(new_n648_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g0493(.A1(new_n678_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g0494(.A1(new_n559_), .A2(new_n560_), .ZN(new_n687_));
  AOI21_X1  g0495(.A(KEYINPUT24), .B1(new_n687_), .B2(new_n531_), .ZN(new_n688_));
  OAI21_X1  g0496(.A(new_n647_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g0497(.A1(new_n452_), .A2(new_n258_), .ZN(new_n690_));
  INV_X1    g0498(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g0499(.A1(new_n556_), .A2(new_n646_), .ZN(new_n692_));
  INV_X1    g0500(.A(KEYINPUT24), .ZN(new_n693_));
  NAND2_X1  g0501(.A1(new_n556_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g0502(.A1(new_n692_), .A2(new_n694_), .A3(new_n678_), .A4(new_n685_), .ZN(new_n695_));
  AND3_X1   g0503(.A1(new_n689_), .A2(new_n691_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g0504(.A(new_n691_), .B1(new_n689_), .B2(new_n695_), .ZN(new_n697_));
  OAI21_X1  g0505(.A(new_n645_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g0506(.A1(new_n689_), .A2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g0507(.A1(new_n699_), .A2(new_n690_), .ZN(new_n700_));
  NAND2_X1  g0508(.A1(new_n573_), .A2(new_n568_), .ZN(new_n701_));
  NAND3_X1  g0509(.A1(new_n689_), .A2(new_n691_), .A3(new_n695_), .ZN(new_n702_));
  NAND3_X1  g0510(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NOR2_X1   g0511(.A1(new_n300_), .A2(new_n310_), .ZN(new_n704_));
  NAND3_X1  g0512(.A1(new_n698_), .A2(new_n703_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g0513(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g0514(.A(new_n704_), .B1(new_n698_), .B2(new_n703_), .ZN(new_n707_));
  NOR2_X1   g0515(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g0516(.A(new_n483_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n709_));
  AOI21_X1  g0517(.A(new_n576_), .B1(new_n709_), .B2(new_n482_), .ZN(new_n710_));
  INV_X1    g0518(.A(KEYINPUT23), .ZN(new_n711_));
  AOI21_X1  g0519(.A(new_n574_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g0520(.A(KEYINPUT23), .B1(new_n575_), .B2(new_n576_), .ZN(new_n713_));
  AOI22_X1  g0521(.A1(new_n580_), .A2(new_n582_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g0522(.A(KEYINPUT27), .ZN(new_n715_));
  NOR2_X1   g0523(.A1(new_n707_), .A2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g0524(.A(new_n708_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  NOR3_X1   g0525(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n718_));
  AOI22_X1  g0526(.A1(new_n485_), .A2(new_n578_), .B1(new_n573_), .B2(new_n571_), .ZN(new_n719_));
  OAI21_X1  g0527(.A(new_n582_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g0528(.A1(new_n712_), .A2(new_n713_), .ZN(new_n721_));
  NAND2_X1  g0529(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g0530(.A1(new_n698_), .A2(new_n703_), .ZN(new_n723_));
  INV_X1    g0531(.A(new_n704_), .ZN(new_n724_));
  NAND2_X1  g0532(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g0533(.A1(new_n725_), .A2(KEYINPUT27), .ZN(new_n726_));
  NAND2_X1  g0534(.A1(new_n725_), .A2(new_n705_), .ZN(new_n727_));
  NAND3_X1  g0535(.A1(new_n722_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g0536(.A(new_n643_), .B1(new_n717_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g0537(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g0538(.A1(new_n717_), .A2(new_n728_), .A3(new_n643_), .ZN(new_n731_));
  NAND2_X1  g0539(.A1(new_n588_), .A2(KEYINPUT22), .ZN(new_n732_));
  NAND3_X1  g0540(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g0541(.A1(new_n592_), .A2(new_n588_), .ZN(new_n734_));
  INV_X1    g0542(.A(new_n734_), .ZN(new_n735_));
  NAND2_X1  g0543(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g0544(.A1(new_n215_), .A2(new_n601_), .ZN(new_n737_));
  INV_X1    g0545(.A(new_n737_), .ZN(new_n738_));
  AND3_X1   g0546(.A1(new_n717_), .A2(new_n728_), .A3(new_n643_), .ZN(new_n739_));
  NOR2_X1   g0547(.A1(new_n739_), .A2(new_n729_), .ZN(new_n740_));
  NAND3_X1  g0548(.A1(new_n740_), .A2(new_n734_), .A3(new_n732_), .ZN(new_n741_));
  NAND3_X1  g0549(.A1(new_n736_), .A2(new_n738_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g0550(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g0551(.A(new_n738_), .B1(new_n736_), .B2(new_n741_), .ZN(new_n744_));
  OAI22_X1  g0552(.A1(new_n640_), .A2(new_n641_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI22_X1  g0553(.A1(new_n638_), .A2(KEYINPUT21), .B1(new_n600_), .B2(new_n603_), .ZN(new_n746_));
  NAND2_X1  g0554(.A1(new_n736_), .A2(new_n741_), .ZN(new_n747_));
  NAND2_X1  g0555(.A1(new_n747_), .A2(new_n737_), .ZN(new_n748_));
  INV_X1    g0556(.A(KEYINPUT21), .ZN(new_n749_));
  NAND4_X1  g0557(.A1(new_n636_), .A2(new_n637_), .A3(new_n749_), .A4(new_n529_), .ZN(new_n750_));
  NAND4_X1  g0558(.A1(new_n746_), .A2(new_n748_), .A3(new_n742_), .A4(new_n750_), .ZN(new_n751_));
  AOI21_X1  g0559(.A(new_n634_), .B1(new_n745_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g0560(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g0561(.A1(new_n745_), .A2(new_n634_), .A3(new_n751_), .ZN(new_n754_));
  NAND2_X1  g0562(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g0563(.A1(new_n631_), .A2(new_n633_), .A3(new_n755_), .ZN(new_n756_));
  AND2_X1   g0564(.A1(new_n632_), .A2(new_n616_), .ZN(new_n757_));
  OAI211_X1 g0565(.A(new_n753_), .B(new_n754_), .C1(new_n757_), .C2(new_n619_), .ZN(new_n758_));
  NAND2_X1  g0566(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g0567(.A1(new_n759_), .A2(G18gat), .A3(G426gat), .ZN(new_n760_));
  NAND2_X1  g0568(.A1(G18gat), .A2(G426gat), .ZN(new_n761_));
  NAND3_X1  g0569(.A1(new_n756_), .A2(new_n758_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g0570(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g0571(.A1(new_n630_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g0572(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g0573(.A1(new_n630_), .A2(new_n763_), .ZN(new_n766_));
  NOR2_X1   g0574(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g0575(.A(G443gat), .ZN(new_n768_));
  NOR2_X1   g0576(.A1(new_n193_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g0577(.A(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g0578(.A(new_n767_), .B(new_n770_), .ZN(G4591gat));
  INV_X1    g0579(.A(KEYINPUT30), .ZN(new_n772_));
  NAND2_X1  g0580(.A1(new_n755_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g0581(.A1(new_n753_), .A2(KEYINPUT30), .A3(new_n754_), .ZN(new_n774_));
  OAI211_X1 g0582(.A(new_n773_), .B(new_n774_), .C1(new_n619_), .C2(new_n757_), .ZN(new_n775_));
  AND2_X1   g0583(.A1(new_n762_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g0584(.A1(new_n205_), .A2(new_n624_), .ZN(new_n777_));
  INV_X1    g0585(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g0586(.A1(new_n753_), .A2(KEYINPUT37), .ZN(new_n779_));
  NOR2_X1   g0587(.A1(new_n640_), .A2(new_n641_), .ZN(new_n780_));
  NOR3_X1   g0588(.A1(new_n780_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n781_));
  INV_X1    g0589(.A(KEYINPUT37), .ZN(new_n782_));
  AOI21_X1  g0590(.A(new_n781_), .B1(new_n752_), .B2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g0591(.A1(new_n215_), .A2(new_n613_), .ZN(new_n784_));
  INV_X1    g0592(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g0593(.A1(new_n740_), .A2(new_n734_), .ZN(new_n786_));
  NAND2_X1  g0594(.A1(new_n742_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g0595(.A1(new_n722_), .A2(new_n727_), .ZN(new_n788_));
  NAND3_X1  g0596(.A1(new_n692_), .A2(new_n678_), .A3(new_n685_), .ZN(new_n789_));
  NAND2_X1  g0597(.A1(new_n702_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g0598(.A(KEYINPUT33), .ZN(new_n791_));
  NAND2_X1  g0599(.A1(new_n680_), .A2(new_n682_), .ZN(new_n792_));
  NAND2_X1  g0600(.A1(new_n792_), .A2(new_n676_), .ZN(new_n793_));
  NOR2_X1   g0601(.A1(new_n651_), .A2(new_n232_), .ZN(new_n794_));
  NAND2_X1  g0602(.A1(G154gat), .A2(G307gat), .ZN(new_n795_));
  INV_X1    g0603(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g0604(.A1(new_n796_), .A2(KEYINPUT32), .ZN(new_n797_));
  NAND2_X1  g0605(.A1(G188gat), .A2(G273gat), .ZN(new_n798_));
  INV_X1    g0606(.A(G171gat), .ZN(new_n799_));
  OAI21_X1  g0607(.A(new_n798_), .B1(new_n799_), .B2(new_n198_), .ZN(new_n800_));
  NAND4_X1  g0608(.A1(G171gat), .A2(G188gat), .A3(G273gat), .A4(G290gat), .ZN(new_n801_));
  AOI21_X1  g0609(.A(new_n661_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AND4_X1   g0610(.A1(G171gat), .A2(G188gat), .A3(G273gat), .A4(G290gat), .ZN(new_n803_));
  NOR2_X1   g0611(.A1(new_n803_), .A2(new_n657_), .ZN(new_n804_));
  OAI21_X1  g0612(.A(new_n797_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g0613(.A1(new_n656_), .A2(new_n657_), .ZN(new_n806_));
  AOI22_X1  g0614(.A1(new_n653_), .A2(new_n666_), .B1(new_n806_), .B2(new_n537_), .ZN(new_n807_));
  AOI22_X1  g0615(.A1(G171gat), .A2(G290gat), .B1(G188gat), .B2(G273gat), .ZN(new_n808_));
  OAI21_X1  g0616(.A(new_n657_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g0617(.A1(new_n661_), .A2(new_n801_), .ZN(new_n810_));
  INV_X1    g0618(.A(KEYINPUT32), .ZN(new_n811_));
  XNOR2_X1  g0619(.A(new_n795_), .B(new_n811_), .ZN(new_n812_));
  NAND3_X1  g0620(.A1(new_n809_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  AND3_X1   g0621(.A1(new_n805_), .A2(new_n807_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g0622(.A(new_n807_), .B1(new_n805_), .B2(new_n813_), .ZN(new_n815_));
  OAI21_X1  g0623(.A(new_n794_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g0624(.A(new_n807_), .ZN(new_n817_));
  INV_X1    g0625(.A(new_n813_), .ZN(new_n818_));
  AOI22_X1  g0626(.A1(new_n809_), .A2(new_n810_), .B1(KEYINPUT32), .B2(new_n796_), .ZN(new_n819_));
  OAI21_X1  g0627(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g0628(.A(new_n794_), .ZN(new_n821_));
  NAND3_X1  g0629(.A1(new_n805_), .A2(new_n807_), .A3(new_n813_), .ZN(new_n822_));
  NAND3_X1  g0630(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g0631(.A1(new_n816_), .A2(new_n823_), .ZN(new_n824_));
  AND3_X1   g0632(.A1(new_n678_), .A2(new_n793_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g0633(.A(new_n824_), .B1(new_n678_), .B2(new_n793_), .ZN(new_n826_));
  OAI21_X1  g0634(.A(new_n791_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g0635(.A1(new_n532_), .A2(new_n258_), .ZN(new_n828_));
  NOR3_X1   g0636(.A1(new_n814_), .A2(new_n815_), .A3(new_n794_), .ZN(new_n829_));
  AOI21_X1  g0637(.A(new_n821_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n830_));
  NOR2_X1   g0638(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g0639(.A(new_n648_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n832_));
  AND2_X1   g0640(.A1(new_n792_), .A2(new_n676_), .ZN(new_n833_));
  OAI21_X1  g0641(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g0642(.A1(new_n678_), .A2(new_n824_), .A3(new_n793_), .ZN(new_n835_));
  NAND3_X1  g0643(.A1(new_n834_), .A2(KEYINPUT33), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g0644(.A1(new_n827_), .A2(new_n828_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g0645(.A(new_n828_), .ZN(new_n838_));
  NAND3_X1  g0646(.A1(new_n834_), .A2(new_n838_), .A3(new_n835_), .ZN(new_n839_));
  NAND3_X1  g0647(.A1(new_n790_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g0648(.A1(new_n299_), .A2(G103gat), .ZN(new_n841_));
  INV_X1    g0649(.A(new_n839_), .ZN(new_n842_));
  AOI21_X1  g0650(.A(new_n838_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n843_));
  OAI211_X1 g0651(.A(new_n702_), .B(new_n789_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  AND3_X1   g0652(.A1(new_n840_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g0653(.A(new_n841_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n846_));
  OAI21_X1  g0654(.A(KEYINPUT34), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g0655(.A1(new_n698_), .A2(new_n703_), .A3(new_n724_), .ZN(new_n848_));
  INV_X1    g0656(.A(KEYINPUT31), .ZN(new_n849_));
  NAND2_X1  g0657(.A1(new_n703_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g0658(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT31), .A4(new_n702_), .ZN(new_n851_));
  NAND3_X1  g0659(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g0660(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g0661(.A1(new_n840_), .A2(new_n844_), .ZN(new_n854_));
  INV_X1    g0662(.A(KEYINPUT34), .ZN(new_n855_));
  NAND3_X1  g0663(.A1(new_n854_), .A2(new_n855_), .A3(new_n841_), .ZN(new_n856_));
  NAND3_X1  g0664(.A1(new_n847_), .A2(new_n853_), .A3(new_n856_), .ZN(new_n857_));
  NOR2_X1   g0665(.A1(new_n310_), .A2(new_n355_), .ZN(new_n858_));
  OAI21_X1  g0666(.A(new_n852_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n859_));
  AND3_X1   g0667(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g0668(.A(new_n858_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n861_));
  OAI211_X1 g0669(.A(new_n731_), .B(new_n788_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g0670(.A1(new_n731_), .A2(new_n788_), .ZN(new_n863_));
  NAND2_X1  g0671(.A1(new_n857_), .A2(new_n859_), .ZN(new_n864_));
  INV_X1    g0672(.A(new_n858_), .ZN(new_n865_));
  NAND2_X1  g0673(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g0674(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n867_));
  NAND3_X1  g0675(.A1(new_n863_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g0676(.A1(new_n862_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g0677(.A1(new_n241_), .A2(new_n601_), .ZN(new_n870_));
  NAND2_X1  g0678(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g0679(.A(new_n870_), .ZN(new_n872_));
  NAND3_X1  g0680(.A1(new_n862_), .A2(new_n868_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g0681(.A(KEYINPUT35), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g0682(.A1(new_n862_), .A2(new_n868_), .A3(KEYINPUT35), .ZN(new_n875_));
  INV_X1    g0683(.A(new_n875_), .ZN(new_n876_));
  OAI211_X1 g0684(.A(new_n787_), .B(KEYINPUT36), .C1(new_n874_), .C2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g0685(.A1(new_n871_), .A2(new_n873_), .ZN(new_n878_));
  NOR2_X1   g0686(.A1(new_n787_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g0687(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g0688(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g0689(.A(KEYINPUT35), .ZN(new_n882_));
  AND3_X1   g0690(.A1(new_n862_), .A2(new_n868_), .A3(new_n872_), .ZN(new_n883_));
  AOI21_X1  g0691(.A(new_n872_), .B1(new_n862_), .B2(new_n868_), .ZN(new_n884_));
  OAI21_X1  g0692(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI22_X1  g0693(.A1(new_n885_), .A2(new_n875_), .B1(new_n742_), .B2(new_n786_), .ZN(new_n886_));
  NOR2_X1   g0694(.A1(new_n886_), .A2(KEYINPUT36), .ZN(new_n887_));
  OAI21_X1  g0695(.A(new_n785_), .B1(new_n881_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g0696(.A(new_n879_), .B1(new_n886_), .B2(KEYINPUT36), .ZN(new_n889_));
  OAI21_X1  g0697(.A(new_n787_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n890_));
  INV_X1    g0698(.A(KEYINPUT36), .ZN(new_n891_));
  NAND2_X1  g0699(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g0700(.A1(new_n889_), .A2(new_n784_), .A3(new_n892_), .ZN(new_n893_));
  AOI22_X1  g0701(.A1(new_n779_), .A2(new_n783_), .B1(new_n888_), .B2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g0702(.A1(new_n752_), .A2(new_n781_), .ZN(new_n895_));
  AND3_X1   g0703(.A1(new_n888_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  OAI21_X1  g0704(.A(new_n778_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g0705(.A1(new_n779_), .A2(new_n783_), .ZN(new_n898_));
  NAND2_X1  g0706(.A1(new_n888_), .A2(new_n893_), .ZN(new_n899_));
  NAND2_X1  g0707(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g0708(.A1(new_n888_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n901_));
  NAND3_X1  g0709(.A1(new_n900_), .A2(new_n777_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g0710(.A1(new_n897_), .A2(new_n902_), .ZN(new_n903_));
  AND2_X1   g0711(.A1(new_n776_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g0712(.A1(new_n776_), .A2(new_n903_), .ZN(new_n905_));
  NOR2_X1   g0713(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g0714(.A1(new_n196_), .A2(new_n768_), .ZN(new_n907_));
  NOR2_X1   g0715(.A1(new_n907_), .A2(KEYINPUT38), .ZN(new_n908_));
  INV_X1    g0716(.A(new_n908_), .ZN(new_n909_));
  NAND2_X1  g0717(.A1(new_n906_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g0718(.A(new_n766_), .B1(new_n770_), .B2(new_n764_), .ZN(new_n911_));
  AND2_X1   g0719(.A1(new_n907_), .A2(KEYINPUT38), .ZN(new_n912_));
  OAI22_X1  g0720(.A1(new_n905_), .A2(new_n904_), .B1(new_n908_), .B2(new_n912_), .ZN(new_n913_));
  NAND3_X1  g0721(.A1(new_n910_), .A2(new_n911_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g0722(.A(new_n914_), .ZN(new_n915_));
  AOI21_X1  g0723(.A(new_n911_), .B1(new_n910_), .B2(new_n913_), .ZN(new_n916_));
  NOR2_X1   g0724(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g0725(.A(G460gat), .ZN(new_n918_));
  NOR2_X1   g0726(.A1(new_n193_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g0727(.A(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g0728(.A(new_n917_), .B(new_n920_), .ZN(G4946gat));
  NAND2_X1  g0729(.A1(G1gat), .A2(G477gat), .ZN(new_n922_));
  XOR2_X1   g0730(.A(new_n922_), .B(KEYINPUT43), .Z(new_n923_));
  INV_X1    g0731(.A(new_n923_), .ZN(new_n924_));
  NAND2_X1  g0732(.A1(new_n776_), .A2(new_n903_), .ZN(new_n925_));
  INV_X1    g0733(.A(new_n907_), .ZN(new_n926_));
  AOI21_X1  g0734(.A(new_n905_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g0735(.A1(new_n205_), .A2(new_n768_), .ZN(new_n928_));
  INV_X1    g0736(.A(new_n928_), .ZN(new_n929_));
  NAND2_X1  g0737(.A1(new_n875_), .A2(new_n872_), .ZN(new_n930_));
  AOI21_X1  g0738(.A(KEYINPUT35), .B1(new_n862_), .B2(new_n868_), .ZN(new_n931_));
  OAI21_X1  g0739(.A(KEYINPUT39), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g0740(.A1(new_n840_), .A2(new_n841_), .A3(new_n844_), .ZN(new_n933_));
  NOR2_X1   g0741(.A1(new_n842_), .A2(new_n843_), .ZN(new_n934_));
  NAND2_X1  g0742(.A1(new_n934_), .A2(new_n790_), .ZN(new_n935_));
  NAND2_X1  g0743(.A1(new_n933_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g0744(.A1(new_n300_), .A2(new_n532_), .ZN(new_n937_));
  AND3_X1   g0745(.A1(new_n834_), .A2(KEYINPUT33), .A3(new_n835_), .ZN(new_n938_));
  AOI21_X1  g0746(.A(KEYINPUT33), .B1(new_n834_), .B2(new_n835_), .ZN(new_n939_));
  OAI21_X1  g0747(.A(new_n838_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  OAI21_X1  g0748(.A(new_n820_), .B1(new_n814_), .B2(new_n794_), .ZN(new_n941_));
  INV_X1    g0749(.A(new_n941_), .ZN(new_n942_));
  NAND2_X1  g0750(.A1(G188gat), .A2(G290gat), .ZN(new_n943_));
  INV_X1    g0751(.A(G205gat), .ZN(new_n944_));
  OAI21_X1  g0752(.A(new_n943_), .B1(new_n944_), .B2(new_n194_), .ZN(new_n945_));
  NAND4_X1  g0753(.A1(G188gat), .A2(G205gat), .A3(G273gat), .A4(G290gat), .ZN(new_n946_));
  NAND2_X1  g0754(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g0755(.A1(new_n947_), .A2(new_n801_), .ZN(new_n948_));
  NOR2_X1   g0756(.A1(new_n799_), .A2(new_n211_), .ZN(new_n949_));
  INV_X1    g0757(.A(new_n949_), .ZN(new_n950_));
  NAND2_X1  g0758(.A1(new_n803_), .A2(new_n946_), .ZN(new_n951_));
  NAND3_X1  g0759(.A1(new_n948_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  AOI21_X1  g0760(.A(new_n803_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n953_));
  INV_X1    g0761(.A(new_n946_), .ZN(new_n954_));
  NOR2_X1   g0762(.A1(new_n954_), .A2(new_n801_), .ZN(new_n955_));
  OAI21_X1  g0763(.A(new_n949_), .B1(new_n953_), .B2(new_n955_), .ZN(new_n956_));
  AOI21_X1  g0764(.A(new_n804_), .B1(new_n809_), .B2(new_n796_), .ZN(new_n957_));
  AND3_X1   g0765(.A1(new_n952_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g0766(.A(new_n957_), .B1(new_n952_), .B2(new_n956_), .ZN(new_n959_));
  INV_X1    g0767(.A(G154gat), .ZN(new_n960_));
  NOR2_X1   g0768(.A1(new_n960_), .A2(new_n232_), .ZN(new_n961_));
  NOR3_X1   g0769(.A1(new_n958_), .A2(new_n959_), .A3(new_n961_), .ZN(new_n962_));
  INV_X1    g0770(.A(new_n961_), .ZN(new_n963_));
  NAND2_X1  g0771(.A1(new_n952_), .A2(new_n956_), .ZN(new_n964_));
  INV_X1    g0772(.A(new_n957_), .ZN(new_n965_));
  NAND2_X1  g0773(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NAND3_X1  g0774(.A1(new_n952_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n967_));
  AOI21_X1  g0775(.A(new_n963_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g0776(.A(new_n942_), .B1(new_n962_), .B2(new_n968_), .ZN(new_n969_));
  OAI21_X1  g0777(.A(new_n961_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n970_));
  NAND3_X1  g0778(.A1(new_n966_), .A2(new_n963_), .A3(new_n967_), .ZN(new_n971_));
  NAND3_X1  g0779(.A1(new_n970_), .A2(new_n971_), .A3(new_n941_), .ZN(new_n972_));
  OAI211_X1 g0780(.A(new_n969_), .B(new_n972_), .C1(new_n651_), .C2(new_n258_), .ZN(new_n973_));
  NOR2_X1   g0781(.A1(new_n651_), .A2(new_n258_), .ZN(new_n974_));
  AND3_X1   g0782(.A1(new_n970_), .A2(new_n971_), .A3(new_n941_), .ZN(new_n975_));
  AOI21_X1  g0783(.A(new_n941_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n976_));
  OAI21_X1  g0784(.A(new_n974_), .B1(new_n975_), .B2(new_n976_), .ZN(new_n977_));
  NAND2_X1  g0785(.A1(new_n973_), .A2(new_n977_), .ZN(new_n978_));
  NOR2_X1   g0786(.A1(new_n978_), .A2(new_n826_), .ZN(new_n979_));
  NAND2_X1  g0787(.A1(new_n940_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g0788(.A1(new_n839_), .A2(new_n834_), .ZN(new_n981_));
  NAND2_X1  g0789(.A1(new_n981_), .A2(new_n978_), .ZN(new_n982_));
  AOI21_X1  g0790(.A(new_n937_), .B1(new_n980_), .B2(new_n982_), .ZN(new_n983_));
  INV_X1    g0791(.A(new_n983_), .ZN(new_n984_));
  AOI22_X1  g0792(.A1(new_n940_), .A2(new_n979_), .B1(new_n978_), .B2(new_n981_), .ZN(new_n985_));
  NAND2_X1  g0793(.A1(new_n985_), .A2(new_n937_), .ZN(new_n986_));
  NAND3_X1  g0794(.A1(new_n936_), .A2(new_n984_), .A3(new_n986_), .ZN(new_n987_));
  AND3_X1   g0795(.A1(new_n980_), .A2(new_n937_), .A3(new_n982_), .ZN(new_n988_));
  OAI211_X1 g0796(.A(new_n933_), .B(new_n935_), .C1(new_n988_), .C2(new_n983_), .ZN(new_n989_));
  NAND2_X1  g0797(.A1(new_n987_), .A2(new_n989_), .ZN(new_n990_));
  NOR2_X1   g0798(.A1(new_n452_), .A2(new_n355_), .ZN(new_n991_));
  NAND2_X1  g0799(.A1(new_n990_), .A2(new_n991_), .ZN(new_n992_));
  INV_X1    g0800(.A(new_n991_), .ZN(new_n993_));
  NAND3_X1  g0801(.A1(new_n987_), .A2(new_n989_), .A3(new_n993_), .ZN(new_n994_));
  NAND2_X1  g0802(.A1(new_n992_), .A2(new_n994_), .ZN(new_n995_));
  INV_X1    g0803(.A(KEYINPUT40), .ZN(new_n996_));
  NAND2_X1  g0804(.A1(new_n852_), .A2(new_n996_), .ZN(new_n997_));
  NAND4_X1  g0805(.A1(new_n848_), .A2(KEYINPUT40), .A3(new_n850_), .A4(new_n851_), .ZN(new_n998_));
  NAND2_X1  g0806(.A1(new_n997_), .A2(new_n998_), .ZN(new_n999_));
  NAND2_X1  g0807(.A1(new_n847_), .A2(new_n856_), .ZN(new_n1000_));
  NOR2_X1   g0808(.A1(new_n999_), .A2(new_n1000_), .ZN(new_n1001_));
  INV_X1    g0809(.A(new_n1001_), .ZN(new_n1002_));
  NAND3_X1  g0810(.A1(new_n995_), .A2(new_n866_), .A3(new_n1002_), .ZN(new_n1003_));
  OAI211_X1 g0811(.A(new_n994_), .B(new_n992_), .C1(new_n861_), .C2(new_n1001_), .ZN(new_n1004_));
  NAND2_X1  g0812(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1005_));
  NOR2_X1   g0813(.A1(new_n310_), .A2(new_n601_), .ZN(new_n1006_));
  NAND2_X1  g0814(.A1(new_n1005_), .A2(new_n1006_), .ZN(new_n1007_));
  INV_X1    g0815(.A(new_n1006_), .ZN(new_n1008_));
  NAND3_X1  g0816(.A1(new_n1003_), .A2(new_n1004_), .A3(new_n1008_), .ZN(new_n1009_));
  AND3_X1   g0817(.A1(new_n1007_), .A2(new_n868_), .A3(new_n1009_), .ZN(new_n1010_));
  NAND2_X1  g0818(.A1(new_n869_), .A2(new_n882_), .ZN(new_n1011_));
  INV_X1    g0819(.A(KEYINPUT39), .ZN(new_n1012_));
  NAND4_X1  g0820(.A1(new_n1011_), .A2(new_n1012_), .A3(new_n875_), .A4(new_n872_), .ZN(new_n1013_));
  NAND3_X1  g0821(.A1(new_n932_), .A2(new_n1010_), .A3(new_n1013_), .ZN(new_n1014_));
  NAND2_X1  g0822(.A1(new_n1007_), .A2(new_n1009_), .ZN(new_n1015_));
  NAND2_X1  g0823(.A1(new_n873_), .A2(new_n868_), .ZN(new_n1016_));
  NAND2_X1  g0824(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  NAND2_X1  g0825(.A1(new_n1014_), .A2(new_n1017_), .ZN(new_n1018_));
  NOR2_X1   g0826(.A1(new_n241_), .A2(new_n613_), .ZN(new_n1019_));
  INV_X1    g0827(.A(new_n1019_), .ZN(new_n1020_));
  NAND2_X1  g0828(.A1(new_n1018_), .A2(new_n1020_), .ZN(new_n1021_));
  NAND3_X1  g0829(.A1(new_n1014_), .A2(new_n1019_), .A3(new_n1017_), .ZN(new_n1022_));
  AOI21_X1  g0830(.A(new_n784_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n1023_));
  AOI21_X1  g0831(.A(new_n878_), .B1(new_n742_), .B2(new_n786_), .ZN(new_n1024_));
  OAI211_X1 g0832(.A(new_n1021_), .B(new_n1022_), .C1(new_n1023_), .C2(new_n1024_), .ZN(new_n1025_));
  NAND2_X1  g0833(.A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1026_));
  INV_X1    g0834(.A(new_n1024_), .ZN(new_n1027_));
  NAND3_X1  g0835(.A1(new_n1026_), .A2(new_n888_), .A3(new_n1027_), .ZN(new_n1028_));
  NAND2_X1  g0836(.A1(new_n1025_), .A2(new_n1028_), .ZN(new_n1029_));
  NOR2_X1   g0837(.A1(new_n215_), .A2(new_n624_), .ZN(new_n1030_));
  NAND2_X1  g0838(.A1(new_n1029_), .A2(new_n1030_), .ZN(new_n1031_));
  INV_X1    g0839(.A(new_n1030_), .ZN(new_n1032_));
  NAND3_X1  g0840(.A1(new_n1025_), .A2(new_n1032_), .A3(new_n1028_), .ZN(new_n1033_));
  AOI21_X1  g0841(.A(new_n777_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n1034_));
  AOI21_X1  g0842(.A(new_n899_), .B1(new_n779_), .B2(new_n783_), .ZN(new_n1035_));
  OAI211_X1 g0843(.A(new_n1031_), .B(new_n1033_), .C1(new_n1034_), .C2(new_n1035_), .ZN(new_n1036_));
  INV_X1    g0844(.A(new_n1035_), .ZN(new_n1037_));
  AND3_X1   g0845(.A1(new_n1025_), .A2(new_n1032_), .A3(new_n1028_), .ZN(new_n1038_));
  AOI21_X1  g0846(.A(new_n1032_), .B1(new_n1025_), .B2(new_n1028_), .ZN(new_n1039_));
  OAI211_X1 g0847(.A(new_n897_), .B(new_n1037_), .C1(new_n1038_), .C2(new_n1039_), .ZN(new_n1040_));
  AOI21_X1  g0848(.A(new_n929_), .B1(new_n1036_), .B2(new_n1040_), .ZN(new_n1041_));
  AND3_X1   g0849(.A1(new_n1036_), .A2(new_n1040_), .A3(new_n929_), .ZN(new_n1042_));
  OAI21_X1  g0850(.A(new_n927_), .B1(new_n1041_), .B2(new_n1042_), .ZN(new_n1043_));
  INV_X1    g0851(.A(new_n1043_), .ZN(new_n1044_));
  NOR3_X1   g0852(.A1(new_n927_), .A2(new_n1042_), .A3(new_n1041_), .ZN(new_n1045_));
  NOR2_X1   g0853(.A1(new_n196_), .A2(new_n918_), .ZN(new_n1046_));
  INV_X1    g0854(.A(new_n1046_), .ZN(new_n1047_));
  NOR3_X1   g0855(.A1(new_n1044_), .A2(new_n1045_), .A3(new_n1047_), .ZN(new_n1048_));
  INV_X1    g0856(.A(new_n1041_), .ZN(new_n1049_));
  NAND3_X1  g0857(.A1(new_n1036_), .A2(new_n1040_), .A3(new_n929_), .ZN(new_n1050_));
  NOR2_X1   g0858(.A1(new_n904_), .A2(new_n907_), .ZN(new_n1051_));
  OAI211_X1 g0859(.A(new_n1049_), .B(new_n1050_), .C1(new_n1051_), .C2(new_n905_), .ZN(new_n1052_));
  AOI21_X1  g0860(.A(new_n1046_), .B1(new_n1052_), .B2(new_n1043_), .ZN(new_n1053_));
  OR2_X1    g0861(.A1(new_n1048_), .A2(new_n1053_), .ZN(new_n1054_));
  AOI21_X1  g0862(.A(new_n916_), .B1(new_n920_), .B2(new_n914_), .ZN(new_n1055_));
  NAND3_X1  g0863(.A1(new_n1054_), .A2(KEYINPUT41), .A3(new_n1055_), .ZN(new_n1056_));
  OAI21_X1  g0864(.A(new_n1055_), .B1(new_n1048_), .B2(new_n1053_), .ZN(new_n1057_));
  INV_X1    g0865(.A(KEYINPUT41), .ZN(new_n1058_));
  NAND2_X1  g0866(.A1(new_n1057_), .A2(new_n1058_), .ZN(new_n1059_));
  NAND2_X1  g0867(.A1(new_n1056_), .A2(new_n1059_), .ZN(new_n1060_));
  OR2_X1    g0868(.A1(new_n1048_), .A2(KEYINPUT42), .ZN(new_n1061_));
  NOR2_X1   g0869(.A1(new_n1055_), .A2(new_n1053_), .ZN(new_n1062_));
  NAND2_X1  g0870(.A1(new_n1048_), .A2(KEYINPUT42), .ZN(new_n1063_));
  NAND3_X1  g0871(.A1(new_n1061_), .A2(new_n1062_), .A3(new_n1063_), .ZN(new_n1064_));
  AOI21_X1  g0872(.A(new_n924_), .B1(new_n1060_), .B2(new_n1064_), .ZN(new_n1065_));
  INV_X1    g0873(.A(new_n1065_), .ZN(new_n1066_));
  NAND3_X1  g0874(.A1(new_n1060_), .A2(new_n924_), .A3(new_n1064_), .ZN(new_n1067_));
  NAND2_X1  g0875(.A1(new_n1066_), .A2(new_n1067_), .ZN(G5308gat));
  INV_X1    g0876(.A(new_n1055_), .ZN(new_n1069_));
  NAND2_X1  g0877(.A1(new_n1054_), .A2(new_n1069_), .ZN(new_n1070_));
  NOR2_X1   g0878(.A1(new_n205_), .A2(new_n918_), .ZN(new_n1071_));
  INV_X1    g0879(.A(new_n1071_), .ZN(new_n1072_));
  NOR2_X1   g0880(.A1(new_n215_), .A2(new_n768_), .ZN(new_n1073_));
  AND3_X1   g0881(.A1(new_n987_), .A2(new_n989_), .A3(new_n993_), .ZN(new_n1074_));
  AOI21_X1  g0882(.A(new_n993_), .B1(new_n987_), .B2(new_n989_), .ZN(new_n1075_));
  NOR2_X1   g0883(.A1(new_n1074_), .A2(new_n1075_), .ZN(new_n1076_));
  NOR3_X1   g0884(.A1(new_n1076_), .A2(new_n861_), .A3(new_n1001_), .ZN(new_n1077_));
  OAI21_X1  g0885(.A(new_n1004_), .B1(new_n1077_), .B2(new_n1006_), .ZN(new_n1078_));
  NAND2_X1  g0886(.A1(G103gat), .A2(G392gat), .ZN(new_n1079_));
  AND3_X1   g0887(.A1(new_n936_), .A2(new_n984_), .A3(new_n986_), .ZN(new_n1080_));
  AOI21_X1  g0888(.A(new_n1080_), .B1(new_n993_), .B2(new_n989_), .ZN(new_n1081_));
  AND2_X1   g0889(.A1(new_n973_), .A2(new_n977_), .ZN(new_n1082_));
  NAND2_X1  g0890(.A1(new_n1082_), .A2(new_n981_), .ZN(new_n1083_));
  OAI21_X1  g0891(.A(new_n1083_), .B1(new_n985_), .B2(new_n937_), .ZN(new_n1084_));
  NAND2_X1  g0892(.A1(new_n973_), .A2(new_n972_), .ZN(new_n1085_));
  INV_X1    g0893(.A(new_n1085_), .ZN(new_n1086_));
  INV_X1    g0894(.A(KEYINPUT46), .ZN(new_n1087_));
  NOR2_X1   g0895(.A1(new_n799_), .A2(new_n232_), .ZN(new_n1088_));
  INV_X1    g0896(.A(new_n1088_), .ZN(new_n1089_));
  AND4_X1   g0897(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1090_));
  AOI22_X1  g0898(.A1(G205gat), .A2(G290gat), .B1(G222gat), .B2(G273gat), .ZN(new_n1091_));
  OAI21_X1  g0899(.A(new_n946_), .B1(new_n1090_), .B2(new_n1091_), .ZN(new_n1092_));
  INV_X1    g0900(.A(G188gat), .ZN(new_n1093_));
  NOR2_X1   g0901(.A1(new_n1093_), .A2(new_n211_), .ZN(new_n1094_));
  NAND4_X1  g0902(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1095_));
  NAND2_X1  g0903(.A1(new_n954_), .A2(new_n1095_), .ZN(new_n1096_));
  NAND3_X1  g0904(.A1(new_n1092_), .A2(new_n1094_), .A3(new_n1096_), .ZN(new_n1097_));
  INV_X1    g0905(.A(KEYINPUT45), .ZN(new_n1098_));
  NAND2_X1  g0906(.A1(new_n1092_), .A2(new_n1096_), .ZN(new_n1099_));
  INV_X1    g0907(.A(new_n1094_), .ZN(new_n1100_));
  AOI21_X1  g0908(.A(new_n1098_), .B1(new_n1099_), .B2(new_n1100_), .ZN(new_n1101_));
  AOI211_X1 g0909(.A(KEYINPUT45), .B(new_n1094_), .C1(new_n1092_), .C2(new_n1096_), .ZN(new_n1102_));
  OAI21_X1  g0910(.A(new_n1097_), .B1(new_n1101_), .B2(new_n1102_), .ZN(new_n1103_));
  AOI21_X1  g0911(.A(new_n953_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n1104_));
  INV_X1    g0912(.A(new_n1104_), .ZN(new_n1105_));
  NAND2_X1  g0913(.A1(new_n1103_), .A2(new_n1105_), .ZN(new_n1106_));
  NAND2_X1  g0914(.A1(G205gat), .A2(G290gat), .ZN(new_n1107_));
  NAND2_X1  g0915(.A1(G222gat), .A2(G273gat), .ZN(new_n1108_));
  NAND2_X1  g0916(.A1(new_n1107_), .A2(new_n1108_), .ZN(new_n1109_));
  INV_X1    g0917(.A(new_n798_), .ZN(new_n1110_));
  AND2_X1   g0918(.A1(G205gat), .A2(G290gat), .ZN(new_n1111_));
  AOI22_X1  g0919(.A1(new_n1109_), .A2(new_n1095_), .B1(new_n1110_), .B2(new_n1111_), .ZN(new_n1112_));
  NOR2_X1   g0920(.A1(new_n1090_), .A2(new_n946_), .ZN(new_n1113_));
  OAI21_X1  g0921(.A(new_n1100_), .B1(new_n1112_), .B2(new_n1113_), .ZN(new_n1114_));
  NAND3_X1  g0922(.A1(new_n1104_), .A2(new_n1097_), .A3(new_n1114_), .ZN(new_n1115_));
  AOI21_X1  g0923(.A(new_n1089_), .B1(new_n1106_), .B2(new_n1115_), .ZN(new_n1116_));
  INV_X1    g0924(.A(new_n1097_), .ZN(new_n1117_));
  NAND2_X1  g0925(.A1(new_n1114_), .A2(KEYINPUT45), .ZN(new_n1118_));
  NAND3_X1  g0926(.A1(new_n1099_), .A2(new_n1098_), .A3(new_n1100_), .ZN(new_n1119_));
  AOI21_X1  g0927(.A(new_n1117_), .B1(new_n1118_), .B2(new_n1119_), .ZN(new_n1120_));
  OAI211_X1 g0928(.A(new_n1089_), .B(new_n1115_), .C1(new_n1120_), .C2(new_n1104_), .ZN(new_n1121_));
  INV_X1    g0929(.A(new_n1121_), .ZN(new_n1122_));
  OAI21_X1  g0930(.A(new_n1087_), .B1(new_n1116_), .B2(new_n1122_), .ZN(new_n1123_));
  NOR2_X1   g0931(.A1(new_n962_), .A2(new_n958_), .ZN(new_n1124_));
  INV_X1    g0932(.A(new_n1124_), .ZN(new_n1125_));
  OAI21_X1  g0933(.A(new_n1115_), .B1(new_n1120_), .B2(new_n1104_), .ZN(new_n1126_));
  NAND2_X1  g0934(.A1(new_n1126_), .A2(new_n1088_), .ZN(new_n1127_));
  NAND3_X1  g0935(.A1(new_n1127_), .A2(KEYINPUT46), .A3(new_n1121_), .ZN(new_n1128_));
  NAND3_X1  g0936(.A1(new_n1123_), .A2(new_n1125_), .A3(new_n1128_), .ZN(new_n1129_));
  NOR2_X1   g0937(.A1(new_n960_), .A2(new_n258_), .ZN(new_n1130_));
  INV_X1    g0938(.A(new_n1130_), .ZN(new_n1131_));
  OAI211_X1 g0939(.A(new_n1087_), .B(new_n1124_), .C1(new_n1116_), .C2(new_n1122_), .ZN(new_n1132_));
  AND3_X1   g0940(.A1(new_n1129_), .A2(new_n1131_), .A3(new_n1132_), .ZN(new_n1133_));
  AOI21_X1  g0941(.A(new_n1131_), .B1(new_n1129_), .B2(new_n1132_), .ZN(new_n1134_));
  OAI21_X1  g0942(.A(new_n1086_), .B1(new_n1133_), .B2(new_n1134_), .ZN(new_n1135_));
  NAND2_X1  g0943(.A1(new_n1129_), .A2(new_n1132_), .ZN(new_n1136_));
  NAND2_X1  g0944(.A1(new_n1136_), .A2(new_n1130_), .ZN(new_n1137_));
  NAND3_X1  g0945(.A1(new_n1129_), .A2(new_n1131_), .A3(new_n1132_), .ZN(new_n1138_));
  NAND3_X1  g0946(.A1(new_n1137_), .A2(new_n1085_), .A3(new_n1138_), .ZN(new_n1139_));
  NOR2_X1   g0947(.A1(new_n300_), .A2(new_n651_), .ZN(new_n1140_));
  INV_X1    g0948(.A(new_n1140_), .ZN(new_n1141_));
  AND3_X1   g0949(.A1(new_n1135_), .A2(new_n1139_), .A3(new_n1141_), .ZN(new_n1142_));
  AOI21_X1  g0950(.A(new_n1141_), .B1(new_n1135_), .B2(new_n1139_), .ZN(new_n1143_));
  OAI21_X1  g0951(.A(new_n1084_), .B1(new_n1142_), .B2(new_n1143_), .ZN(new_n1144_));
  NOR3_X1   g0952(.A1(new_n1133_), .A2(new_n1134_), .A3(new_n1086_), .ZN(new_n1145_));
  AOI21_X1  g0953(.A(new_n1085_), .B1(new_n1137_), .B2(new_n1138_), .ZN(new_n1146_));
  OAI21_X1  g0954(.A(new_n1140_), .B1(new_n1145_), .B2(new_n1146_), .ZN(new_n1147_));
  NAND2_X1  g0955(.A1(new_n1082_), .A2(new_n834_), .ZN(new_n1148_));
  AOI21_X1  g0956(.A(new_n828_), .B1(new_n827_), .B2(new_n836_), .ZN(new_n1149_));
  OAI21_X1  g0957(.A(new_n982_), .B1(new_n1148_), .B2(new_n1149_), .ZN(new_n1150_));
  INV_X1    g0958(.A(new_n937_), .ZN(new_n1151_));
  AOI22_X1  g0959(.A1(new_n1150_), .A2(new_n1151_), .B1(new_n1082_), .B2(new_n981_), .ZN(new_n1152_));
  NAND3_X1  g0960(.A1(new_n1135_), .A2(new_n1139_), .A3(new_n1141_), .ZN(new_n1153_));
  NAND3_X1  g0961(.A1(new_n1147_), .A2(new_n1152_), .A3(new_n1153_), .ZN(new_n1154_));
  NAND2_X1  g0962(.A1(G120gat), .A2(G375gat), .ZN(new_n1155_));
  XOR2_X1   g0963(.A(new_n1155_), .B(KEYINPUT47), .Z(new_n1156_));
  AND3_X1   g0964(.A1(new_n1144_), .A2(new_n1154_), .A3(new_n1156_), .ZN(new_n1157_));
  AOI21_X1  g0965(.A(new_n1156_), .B1(new_n1144_), .B2(new_n1154_), .ZN(new_n1158_));
  OAI21_X1  g0966(.A(new_n1081_), .B1(new_n1157_), .B2(new_n1158_), .ZN(new_n1159_));
  NAND2_X1  g0967(.A1(new_n1144_), .A2(new_n1154_), .ZN(new_n1160_));
  NAND2_X1  g0968(.A1(new_n1160_), .A2(new_n1155_), .ZN(new_n1161_));
  INV_X1    g0969(.A(new_n989_), .ZN(new_n1162_));
  OAI21_X1  g0970(.A(new_n987_), .B1(new_n1162_), .B2(new_n991_), .ZN(new_n1163_));
  NAND3_X1  g0971(.A1(new_n1144_), .A2(new_n1154_), .A3(new_n1156_), .ZN(new_n1164_));
  NAND3_X1  g0972(.A1(new_n1161_), .A2(new_n1163_), .A3(new_n1164_), .ZN(new_n1165_));
  AOI21_X1  g0973(.A(new_n1079_), .B1(new_n1159_), .B2(new_n1165_), .ZN(new_n1166_));
  INV_X1    g0974(.A(new_n1166_), .ZN(new_n1167_));
  NAND3_X1  g0975(.A1(new_n1159_), .A2(new_n1165_), .A3(new_n1079_), .ZN(new_n1168_));
  NAND3_X1  g0976(.A1(new_n1078_), .A2(new_n1167_), .A3(new_n1168_), .ZN(new_n1169_));
  AND3_X1   g0977(.A1(new_n1159_), .A2(new_n1165_), .A3(new_n1079_), .ZN(new_n1170_));
  OAI211_X1 g0978(.A(new_n1009_), .B(new_n1004_), .C1(new_n1170_), .C2(new_n1166_), .ZN(new_n1171_));
  NAND2_X1  g0979(.A1(new_n1169_), .A2(new_n1171_), .ZN(new_n1172_));
  NOR2_X1   g0980(.A1(new_n310_), .A2(new_n613_), .ZN(new_n1173_));
  INV_X1    g0981(.A(new_n1173_), .ZN(new_n1174_));
  NAND2_X1  g0982(.A1(new_n1172_), .A2(new_n1174_), .ZN(new_n1175_));
  NAND3_X1  g0983(.A1(new_n1169_), .A2(new_n1171_), .A3(new_n1173_), .ZN(new_n1176_));
  NAND3_X1  g0984(.A1(new_n1175_), .A2(KEYINPUT48), .A3(new_n1176_), .ZN(new_n1177_));
  AOI21_X1  g0985(.A(new_n1015_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n1178_));
  INV_X1    g0986(.A(new_n1178_), .ZN(new_n1179_));
  INV_X1    g0987(.A(KEYINPUT48), .ZN(new_n1180_));
  NAND3_X1  g0988(.A1(new_n1172_), .A2(new_n1180_), .A3(new_n1174_), .ZN(new_n1181_));
  AND3_X1   g0989(.A1(new_n1177_), .A2(new_n1179_), .A3(new_n1181_), .ZN(new_n1182_));
  INV_X1    g0990(.A(KEYINPUT44), .ZN(new_n1183_));
  INV_X1    g0991(.A(new_n1017_), .ZN(new_n1184_));
  NAND3_X1  g0992(.A1(new_n1007_), .A2(new_n868_), .A3(new_n1009_), .ZN(new_n1185_));
  NAND3_X1  g0993(.A1(new_n1011_), .A2(new_n875_), .A3(new_n872_), .ZN(new_n1186_));
  AOI21_X1  g0994(.A(new_n1185_), .B1(new_n1186_), .B2(KEYINPUT39), .ZN(new_n1187_));
  AOI21_X1  g0995(.A(new_n1184_), .B1(new_n1187_), .B2(new_n1013_), .ZN(new_n1188_));
  OAI21_X1  g0996(.A(new_n1183_), .B1(new_n1188_), .B2(new_n1019_), .ZN(new_n1189_));
  AOI21_X1  g0997(.A(new_n1019_), .B1(new_n1014_), .B2(new_n1017_), .ZN(new_n1190_));
  NAND2_X1  g0998(.A1(new_n1190_), .A2(KEYINPUT44), .ZN(new_n1191_));
  NAND3_X1  g0999(.A1(new_n1182_), .A2(new_n1189_), .A3(new_n1191_), .ZN(new_n1192_));
  AND2_X1   g1000(.A1(new_n1175_), .A2(new_n1176_), .ZN(new_n1193_));
  OAI21_X1  g1001(.A(new_n1193_), .B1(new_n1190_), .B2(new_n1178_), .ZN(new_n1194_));
  INV_X1    g1002(.A(KEYINPUT49), .ZN(new_n1195_));
  NAND2_X1  g1003(.A1(new_n1194_), .A2(new_n1195_), .ZN(new_n1196_));
  OAI211_X1 g1004(.A(KEYINPUT49), .B(new_n1193_), .C1(new_n1190_), .C2(new_n1178_), .ZN(new_n1197_));
  NAND3_X1  g1005(.A1(new_n1192_), .A2(new_n1196_), .A3(new_n1197_), .ZN(new_n1198_));
  NOR2_X1   g1006(.A1(new_n241_), .A2(new_n624_), .ZN(new_n1199_));
  INV_X1    g1007(.A(new_n1199_), .ZN(new_n1200_));
  NAND2_X1  g1008(.A1(new_n1198_), .A2(new_n1200_), .ZN(new_n1201_));
  AND3_X1   g1009(.A1(new_n1026_), .A2(new_n888_), .A3(new_n1027_), .ZN(new_n1202_));
  OAI21_X1  g1010(.A(new_n1025_), .B1(new_n1202_), .B2(new_n1030_), .ZN(new_n1203_));
  NAND4_X1  g1011(.A1(new_n1192_), .A2(new_n1196_), .A3(new_n1199_), .A4(new_n1197_), .ZN(new_n1204_));
  AND3_X1   g1012(.A1(new_n1201_), .A2(new_n1203_), .A3(new_n1204_), .ZN(new_n1205_));
  AOI21_X1  g1013(.A(new_n1203_), .B1(new_n1201_), .B2(new_n1204_), .ZN(new_n1206_));
  OAI21_X1  g1014(.A(new_n1073_), .B1(new_n1205_), .B2(new_n1206_), .ZN(new_n1207_));
  NAND2_X1  g1015(.A1(new_n1201_), .A2(new_n1204_), .ZN(new_n1208_));
  INV_X1    g1016(.A(new_n1203_), .ZN(new_n1209_));
  NAND2_X1  g1017(.A1(new_n1208_), .A2(new_n1209_), .ZN(new_n1210_));
  INV_X1    g1018(.A(new_n1073_), .ZN(new_n1211_));
  NAND3_X1  g1019(.A1(new_n1201_), .A2(new_n1203_), .A3(new_n1204_), .ZN(new_n1212_));
  NAND3_X1  g1020(.A1(new_n1210_), .A2(new_n1211_), .A3(new_n1212_), .ZN(new_n1213_));
  AND4_X1   g1021(.A1(new_n1036_), .A2(new_n1207_), .A3(new_n1213_), .A4(new_n1050_), .ZN(new_n1214_));
  AOI22_X1  g1022(.A1(new_n1213_), .A2(new_n1207_), .B1(new_n1050_), .B2(new_n1036_), .ZN(new_n1215_));
  OAI21_X1  g1023(.A(new_n1072_), .B1(new_n1214_), .B2(new_n1215_), .ZN(new_n1216_));
  INV_X1    g1024(.A(new_n1040_), .ZN(new_n1217_));
  OAI21_X1  g1025(.A(new_n1036_), .B1(new_n1217_), .B2(new_n928_), .ZN(new_n1218_));
  NOR3_X1   g1026(.A1(new_n1205_), .A2(new_n1206_), .A3(new_n1073_), .ZN(new_n1219_));
  AOI21_X1  g1027(.A(new_n1211_), .B1(new_n1210_), .B2(new_n1212_), .ZN(new_n1220_));
  OAI21_X1  g1028(.A(new_n1218_), .B1(new_n1219_), .B2(new_n1220_), .ZN(new_n1221_));
  NAND4_X1  g1029(.A1(new_n1207_), .A2(new_n1213_), .A3(new_n1050_), .A4(new_n1036_), .ZN(new_n1222_));
  NAND3_X1  g1030(.A1(new_n1221_), .A2(new_n1071_), .A3(new_n1222_), .ZN(new_n1223_));
  NAND2_X1  g1031(.A1(new_n1216_), .A2(new_n1223_), .ZN(new_n1224_));
  AOI21_X1  g1032(.A(new_n1045_), .B1(new_n1047_), .B2(new_n1043_), .ZN(new_n1225_));
  NAND2_X1  g1033(.A1(new_n1224_), .A2(new_n1225_), .ZN(new_n1226_));
  OAI21_X1  g1034(.A(new_n1052_), .B1(new_n1044_), .B2(new_n1046_), .ZN(new_n1227_));
  NAND3_X1  g1035(.A1(new_n1227_), .A2(new_n1216_), .A3(new_n1223_), .ZN(new_n1228_));
  NAND2_X1  g1036(.A1(new_n1226_), .A2(new_n1228_), .ZN(new_n1229_));
  NAND3_X1  g1037(.A1(new_n1229_), .A2(G18gat), .A3(G477gat), .ZN(new_n1230_));
  NAND2_X1  g1038(.A1(G18gat), .A2(G477gat), .ZN(new_n1231_));
  NAND3_X1  g1039(.A1(new_n1226_), .A2(new_n1228_), .A3(new_n1231_), .ZN(new_n1232_));
  NAND2_X1  g1040(.A1(new_n1230_), .A2(new_n1232_), .ZN(new_n1233_));
  NAND3_X1  g1041(.A1(new_n1066_), .A2(new_n1070_), .A3(new_n1233_), .ZN(new_n1234_));
  INV_X1    g1042(.A(new_n1070_), .ZN(new_n1235_));
  OAI211_X1 g1043(.A(new_n1232_), .B(new_n1230_), .C1(new_n1065_), .C2(new_n1235_), .ZN(new_n1236_));
  NAND2_X1  g1044(.A1(new_n1234_), .A2(new_n1236_), .ZN(new_n1237_));
  NAND2_X1  g1045(.A1(G1gat), .A2(G494gat), .ZN(new_n1238_));
  XNOR2_X1  g1046(.A(new_n1238_), .B(KEYINPUT50), .ZN(new_n1239_));
  NAND2_X1  g1047(.A1(new_n1237_), .A2(new_n1239_), .ZN(new_n1240_));
  INV_X1    g1048(.A(new_n1239_), .ZN(new_n1241_));
  NAND3_X1  g1049(.A1(new_n1234_), .A2(new_n1236_), .A3(new_n1241_), .ZN(new_n1242_));
  NAND2_X1  g1050(.A1(new_n1240_), .A2(new_n1242_), .ZN(G5672gat));
  NAND4_X1  g1051(.A1(new_n1227_), .A2(KEYINPUT51), .A3(new_n1216_), .A4(new_n1223_), .ZN(new_n1244_));
  INV_X1    g1052(.A(KEYINPUT51), .ZN(new_n1245_));
  NAND2_X1  g1053(.A1(new_n1228_), .A2(new_n1245_), .ZN(new_n1246_));
  NAND3_X1  g1054(.A1(new_n1232_), .A2(new_n1244_), .A3(new_n1246_), .ZN(new_n1247_));
  INV_X1    g1055(.A(new_n1247_), .ZN(new_n1248_));
  AOI21_X1  g1056(.A(new_n1205_), .B1(new_n1210_), .B2(new_n1211_), .ZN(new_n1249_));
  INV_X1    g1057(.A(new_n1156_), .ZN(new_n1250_));
  NAND2_X1  g1058(.A1(new_n1160_), .A2(new_n1250_), .ZN(new_n1251_));
  NAND3_X1  g1059(.A1(new_n1251_), .A2(new_n1163_), .A3(new_n1164_), .ZN(new_n1252_));
  NAND2_X1  g1060(.A1(new_n1168_), .A2(new_n1252_), .ZN(new_n1253_));
  INV_X1    g1061(.A(new_n1253_), .ZN(new_n1254_));
  NAND2_X1  g1062(.A1(new_n1084_), .A2(KEYINPUT53), .ZN(new_n1255_));
  AND3_X1   g1063(.A1(new_n1255_), .A2(new_n1153_), .A3(new_n1147_), .ZN(new_n1256_));
  OR2_X1    g1064(.A1(new_n1084_), .A2(KEYINPUT53), .ZN(new_n1257_));
  NAND2_X1  g1065(.A1(new_n1256_), .A2(new_n1257_), .ZN(new_n1258_));
  NAND2_X1  g1066(.A1(new_n1161_), .A2(new_n1258_), .ZN(new_n1259_));
  NOR2_X1   g1067(.A1(new_n300_), .A2(new_n960_), .ZN(new_n1260_));
  INV_X1    g1068(.A(new_n1260_), .ZN(new_n1261_));
  AOI21_X1  g1069(.A(new_n1112_), .B1(new_n1100_), .B2(new_n1096_), .ZN(new_n1262_));
  INV_X1    g1070(.A(new_n1262_), .ZN(new_n1263_));
  NOR2_X1   g1071(.A1(new_n944_), .A2(new_n211_), .ZN(new_n1264_));
  NAND4_X1  g1072(.A1(G222gat), .A2(G239gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1265_));
  NAND2_X1  g1073(.A1(new_n1090_), .A2(new_n1265_), .ZN(new_n1266_));
  AND2_X1   g1074(.A1(G222gat), .A2(G273gat), .ZN(new_n1267_));
  AND2_X1   g1075(.A1(G239gat), .A2(G290gat), .ZN(new_n1268_));
  NAND2_X1  g1076(.A1(G222gat), .A2(G290gat), .ZN(new_n1269_));
  NAND2_X1  g1077(.A1(G239gat), .A2(G273gat), .ZN(new_n1270_));
  AOI22_X1  g1078(.A1(new_n1267_), .A2(new_n1268_), .B1(new_n1269_), .B2(new_n1270_), .ZN(new_n1271_));
  OAI211_X1 g1079(.A(new_n1264_), .B(new_n1266_), .C1(new_n1271_), .C2(new_n1090_), .ZN(new_n1272_));
  INV_X1    g1080(.A(KEYINPUT57), .ZN(new_n1273_));
  NAND2_X1  g1081(.A1(new_n1272_), .A2(new_n1273_), .ZN(new_n1274_));
  NAND2_X1  g1082(.A1(new_n1269_), .A2(new_n1270_), .ZN(new_n1275_));
  NAND2_X1  g1083(.A1(new_n1275_), .A2(new_n1265_), .ZN(new_n1276_));
  NAND2_X1  g1084(.A1(new_n1276_), .A2(new_n1095_), .ZN(new_n1277_));
  NAND4_X1  g1085(.A1(new_n1277_), .A2(KEYINPUT57), .A3(new_n1264_), .A4(new_n1266_), .ZN(new_n1278_));
  NAND2_X1  g1086(.A1(new_n1274_), .A2(new_n1278_), .ZN(new_n1279_));
  INV_X1    g1087(.A(KEYINPUT56), .ZN(new_n1280_));
  AND2_X1   g1088(.A1(G205gat), .A2(G273gat), .ZN(new_n1281_));
  AND2_X1   g1089(.A1(G222gat), .A2(G290gat), .ZN(new_n1282_));
  AOI22_X1  g1090(.A1(new_n1275_), .A2(new_n1265_), .B1(new_n1281_), .B2(new_n1282_), .ZN(new_n1283_));
  AND4_X1   g1091(.A1(G222gat), .A2(G239gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1284_));
  NOR2_X1   g1092(.A1(new_n1284_), .A2(new_n1095_), .ZN(new_n1285_));
  OAI21_X1  g1093(.A(new_n1280_), .B1(new_n1283_), .B2(new_n1285_), .ZN(new_n1286_));
  NAND3_X1  g1094(.A1(new_n1271_), .A2(KEYINPUT56), .A3(new_n1095_), .ZN(new_n1287_));
  AOI21_X1  g1095(.A(new_n1264_), .B1(new_n1286_), .B2(new_n1287_), .ZN(new_n1288_));
  OAI21_X1  g1096(.A(new_n1263_), .B1(new_n1279_), .B2(new_n1288_), .ZN(new_n1289_));
  INV_X1    g1097(.A(new_n1264_), .ZN(new_n1290_));
  AOI21_X1  g1098(.A(KEYINPUT56), .B1(new_n1277_), .B2(new_n1266_), .ZN(new_n1291_));
  INV_X1    g1099(.A(new_n1287_), .ZN(new_n1292_));
  OAI21_X1  g1100(.A(new_n1290_), .B1(new_n1291_), .B2(new_n1292_), .ZN(new_n1293_));
  NAND3_X1  g1101(.A1(new_n1286_), .A2(new_n1264_), .A3(new_n1287_), .ZN(new_n1294_));
  NAND3_X1  g1102(.A1(new_n1293_), .A2(new_n1262_), .A3(new_n1294_), .ZN(new_n1295_));
  NAND2_X1  g1103(.A1(new_n1289_), .A2(new_n1295_), .ZN(new_n1296_));
  NOR2_X1   g1104(.A1(new_n1093_), .A2(new_n232_), .ZN(new_n1297_));
  NAND2_X1  g1105(.A1(new_n1296_), .A2(new_n1297_), .ZN(new_n1298_));
  INV_X1    g1106(.A(new_n1297_), .ZN(new_n1299_));
  NAND3_X1  g1107(.A1(new_n1289_), .A2(new_n1295_), .A3(new_n1299_), .ZN(new_n1300_));
  NAND2_X1  g1108(.A1(new_n1106_), .A2(KEYINPUT55), .ZN(new_n1301_));
  NAND3_X1  g1109(.A1(new_n1298_), .A2(new_n1300_), .A3(new_n1301_), .ZN(new_n1302_));
  NAND2_X1  g1110(.A1(new_n1121_), .A2(new_n1106_), .ZN(new_n1303_));
  INV_X1    g1111(.A(new_n1303_), .ZN(new_n1304_));
  NAND2_X1  g1112(.A1(new_n1302_), .A2(new_n1304_), .ZN(new_n1305_));
  NOR2_X1   g1113(.A1(new_n799_), .A2(new_n258_), .ZN(new_n1306_));
  INV_X1    g1114(.A(new_n1306_), .ZN(new_n1307_));
  NAND4_X1  g1115(.A1(new_n1298_), .A2(new_n1303_), .A3(new_n1300_), .A4(new_n1301_), .ZN(new_n1308_));
  AND3_X1   g1116(.A1(new_n1305_), .A2(new_n1307_), .A3(new_n1308_), .ZN(new_n1309_));
  AOI21_X1  g1117(.A(new_n1307_), .B1(new_n1305_), .B2(new_n1308_), .ZN(new_n1310_));
  NOR2_X1   g1118(.A1(new_n1309_), .A2(new_n1310_), .ZN(new_n1311_));
  NAND3_X1  g1119(.A1(new_n1125_), .A2(new_n1121_), .A3(new_n1127_), .ZN(new_n1312_));
  NAND2_X1  g1120(.A1(new_n1138_), .A2(new_n1312_), .ZN(new_n1313_));
  INV_X1    g1121(.A(KEYINPUT54), .ZN(new_n1314_));
  NAND2_X1  g1122(.A1(new_n1138_), .A2(new_n1314_), .ZN(new_n1315_));
  AND3_X1   g1123(.A1(new_n1311_), .A2(new_n1313_), .A3(new_n1315_), .ZN(new_n1316_));
  AOI21_X1  g1124(.A(new_n1313_), .B1(new_n1311_), .B2(new_n1315_), .ZN(new_n1317_));
  OAI21_X1  g1125(.A(new_n1261_), .B1(new_n1316_), .B2(new_n1317_), .ZN(new_n1318_));
  INV_X1    g1126(.A(new_n1300_), .ZN(new_n1319_));
  AOI21_X1  g1127(.A(new_n1299_), .B1(new_n1289_), .B2(new_n1295_), .ZN(new_n1320_));
  NOR2_X1   g1128(.A1(new_n1319_), .A2(new_n1320_), .ZN(new_n1321_));
  AOI21_X1  g1129(.A(new_n1303_), .B1(new_n1321_), .B2(new_n1301_), .ZN(new_n1322_));
  INV_X1    g1130(.A(new_n1308_), .ZN(new_n1323_));
  OAI21_X1  g1131(.A(new_n1306_), .B1(new_n1322_), .B2(new_n1323_), .ZN(new_n1324_));
  NAND3_X1  g1132(.A1(new_n1305_), .A2(new_n1307_), .A3(new_n1308_), .ZN(new_n1325_));
  NAND2_X1  g1133(.A1(new_n1324_), .A2(new_n1325_), .ZN(new_n1326_));
  OAI211_X1 g1134(.A(new_n1138_), .B(new_n1312_), .C1(new_n1326_), .C2(new_n1314_), .ZN(new_n1327_));
  NAND3_X1  g1135(.A1(new_n1311_), .A2(new_n1313_), .A3(new_n1315_), .ZN(new_n1328_));
  NAND3_X1  g1136(.A1(new_n1327_), .A2(new_n1260_), .A3(new_n1328_), .ZN(new_n1329_));
  NAND2_X1  g1137(.A1(new_n1318_), .A2(new_n1329_), .ZN(new_n1330_));
  INV_X1    g1138(.A(KEYINPUT58), .ZN(new_n1331_));
  NAND2_X1  g1139(.A1(new_n1318_), .A2(new_n1331_), .ZN(new_n1332_));
  NAND2_X1  g1140(.A1(new_n1153_), .A2(new_n1139_), .ZN(new_n1333_));
  NAND3_X1  g1141(.A1(new_n1330_), .A2(new_n1332_), .A3(new_n1333_), .ZN(new_n1334_));
  NOR2_X1   g1142(.A1(new_n651_), .A2(new_n355_), .ZN(new_n1335_));
  INV_X1    g1143(.A(new_n1335_), .ZN(new_n1336_));
  AOI21_X1  g1144(.A(new_n1145_), .B1(new_n1141_), .B2(new_n1135_), .ZN(new_n1337_));
  OAI211_X1 g1145(.A(new_n1318_), .B(new_n1329_), .C1(new_n1337_), .C2(new_n1331_), .ZN(new_n1338_));
  AND3_X1   g1146(.A1(new_n1334_), .A2(new_n1336_), .A3(new_n1338_), .ZN(new_n1339_));
  AOI21_X1  g1147(.A(new_n1336_), .B1(new_n1334_), .B2(new_n1338_), .ZN(new_n1340_));
  OAI21_X1  g1148(.A(new_n1259_), .B1(new_n1339_), .B2(new_n1340_), .ZN(new_n1341_));
  AND2_X1   g1149(.A1(new_n1318_), .A2(new_n1329_), .ZN(new_n1342_));
  AOI21_X1  g1150(.A(new_n1260_), .B1(new_n1327_), .B2(new_n1328_), .ZN(new_n1343_));
  OAI21_X1  g1151(.A(new_n1333_), .B1(new_n1343_), .B2(KEYINPUT58), .ZN(new_n1344_));
  NOR2_X1   g1152(.A1(new_n1342_), .A2(new_n1344_), .ZN(new_n1345_));
  INV_X1    g1153(.A(new_n1338_), .ZN(new_n1346_));
  OAI21_X1  g1154(.A(new_n1335_), .B1(new_n1345_), .B2(new_n1346_), .ZN(new_n1347_));
  NAND3_X1  g1155(.A1(new_n1334_), .A2(new_n1336_), .A3(new_n1338_), .ZN(new_n1348_));
  AOI21_X1  g1156(.A(new_n1158_), .B1(new_n1257_), .B2(new_n1256_), .ZN(new_n1349_));
  NAND3_X1  g1157(.A1(new_n1347_), .A2(new_n1348_), .A3(new_n1349_), .ZN(new_n1350_));
  NOR2_X1   g1158(.A1(new_n532_), .A2(new_n601_), .ZN(new_n1351_));
  INV_X1    g1159(.A(new_n1351_), .ZN(new_n1352_));
  NAND3_X1  g1160(.A1(new_n1341_), .A2(new_n1350_), .A3(new_n1352_), .ZN(new_n1353_));
  AOI21_X1  g1161(.A(new_n1352_), .B1(new_n1341_), .B2(new_n1350_), .ZN(new_n1354_));
  INV_X1    g1162(.A(KEYINPUT59), .ZN(new_n1355_));
  OAI21_X1  g1163(.A(new_n1353_), .B1(new_n1354_), .B2(new_n1355_), .ZN(new_n1356_));
  AOI211_X1 g1164(.A(KEYINPUT59), .B(new_n1352_), .C1(new_n1341_), .C2(new_n1350_), .ZN(new_n1357_));
  OAI21_X1  g1165(.A(new_n1254_), .B1(new_n1356_), .B2(new_n1357_), .ZN(new_n1358_));
  NAND2_X1  g1166(.A1(new_n1251_), .A2(new_n1258_), .ZN(new_n1359_));
  NOR3_X1   g1167(.A1(new_n1339_), .A2(new_n1340_), .A3(new_n1359_), .ZN(new_n1360_));
  AOI22_X1  g1168(.A1(new_n1155_), .A2(new_n1160_), .B1(new_n1256_), .B2(new_n1257_), .ZN(new_n1361_));
  AOI21_X1  g1169(.A(new_n1361_), .B1(new_n1347_), .B2(new_n1348_), .ZN(new_n1362_));
  OAI21_X1  g1170(.A(new_n1351_), .B1(new_n1360_), .B2(new_n1362_), .ZN(new_n1363_));
  NAND3_X1  g1171(.A1(new_n1363_), .A2(new_n1253_), .A3(new_n1353_), .ZN(new_n1364_));
  NAND2_X1  g1172(.A1(new_n1358_), .A2(new_n1364_), .ZN(new_n1365_));
  NOR2_X1   g1173(.A1(new_n452_), .A2(new_n613_), .ZN(new_n1366_));
  NAND2_X1  g1174(.A1(new_n1365_), .A2(new_n1366_), .ZN(new_n1367_));
  INV_X1    g1175(.A(KEYINPUT60), .ZN(new_n1368_));
  INV_X1    g1176(.A(new_n1366_), .ZN(new_n1369_));
  NAND3_X1  g1177(.A1(new_n1358_), .A2(new_n1369_), .A3(new_n1364_), .ZN(new_n1370_));
  NAND3_X1  g1178(.A1(new_n1367_), .A2(new_n1368_), .A3(new_n1370_), .ZN(new_n1371_));
  INV_X1    g1179(.A(new_n1171_), .ZN(new_n1372_));
  OAI21_X1  g1180(.A(new_n1169_), .B1(new_n1372_), .B2(new_n1173_), .ZN(new_n1373_));
  INV_X1    g1181(.A(new_n1373_), .ZN(new_n1374_));
  NAND3_X1  g1182(.A1(new_n1365_), .A2(KEYINPUT60), .A3(new_n1366_), .ZN(new_n1375_));
  NAND3_X1  g1183(.A1(new_n1371_), .A2(new_n1374_), .A3(new_n1375_), .ZN(new_n1376_));
  NOR2_X1   g1184(.A1(new_n310_), .A2(new_n624_), .ZN(new_n1377_));
  NAND3_X1  g1185(.A1(new_n1367_), .A2(new_n1373_), .A3(new_n1370_), .ZN(new_n1378_));
  AND3_X1   g1186(.A1(new_n1376_), .A2(new_n1377_), .A3(new_n1378_), .ZN(new_n1379_));
  AOI21_X1  g1187(.A(new_n1377_), .B1(new_n1376_), .B2(new_n1378_), .ZN(new_n1380_));
  NOR2_X1   g1188(.A1(new_n1379_), .A2(new_n1380_), .ZN(new_n1381_));
  NOR2_X1   g1189(.A1(new_n1190_), .A2(new_n1178_), .ZN(new_n1382_));
  NAND2_X1  g1190(.A1(new_n1177_), .A2(new_n1181_), .ZN(new_n1383_));
  NOR2_X1   g1191(.A1(new_n1382_), .A2(new_n1383_), .ZN(new_n1384_));
  INV_X1    g1192(.A(new_n1384_), .ZN(new_n1385_));
  NAND2_X1  g1193(.A1(new_n1201_), .A2(new_n1385_), .ZN(new_n1386_));
  NAND2_X1  g1194(.A1(new_n1381_), .A2(new_n1386_), .ZN(new_n1387_));
  NOR2_X1   g1195(.A1(new_n241_), .A2(new_n768_), .ZN(new_n1388_));
  INV_X1    g1196(.A(new_n1388_), .ZN(new_n1389_));
  AOI21_X1  g1197(.A(new_n1384_), .B1(new_n1198_), .B2(new_n1200_), .ZN(new_n1390_));
  OAI21_X1  g1198(.A(new_n1390_), .B1(new_n1380_), .B2(new_n1379_), .ZN(new_n1391_));
  AND3_X1   g1199(.A1(new_n1387_), .A2(new_n1389_), .A3(new_n1391_), .ZN(new_n1392_));
  AOI21_X1  g1200(.A(new_n1389_), .B1(new_n1387_), .B2(new_n1391_), .ZN(new_n1393_));
  OAI21_X1  g1201(.A(new_n1249_), .B1(new_n1392_), .B2(new_n1393_), .ZN(new_n1394_));
  NOR2_X1   g1202(.A1(new_n1381_), .A2(new_n1386_), .ZN(new_n1395_));
  NOR3_X1   g1203(.A1(new_n1390_), .A2(new_n1379_), .A3(new_n1380_), .ZN(new_n1396_));
  OAI21_X1  g1204(.A(new_n1388_), .B1(new_n1395_), .B2(new_n1396_), .ZN(new_n1397_));
  OAI21_X1  g1205(.A(new_n1212_), .B1(new_n1206_), .B2(new_n1073_), .ZN(new_n1398_));
  NAND3_X1  g1206(.A1(new_n1387_), .A2(new_n1389_), .A3(new_n1391_), .ZN(new_n1399_));
  NAND3_X1  g1207(.A1(new_n1397_), .A2(new_n1398_), .A3(new_n1399_), .ZN(new_n1400_));
  NOR2_X1   g1208(.A1(new_n215_), .A2(new_n918_), .ZN(new_n1401_));
  AND3_X1   g1209(.A1(new_n1394_), .A2(new_n1400_), .A3(new_n1401_), .ZN(new_n1402_));
  XOR2_X1   g1210(.A(new_n1401_), .B(KEYINPUT61), .Z(new_n1403_));
  AOI21_X1  g1211(.A(new_n1403_), .B1(new_n1394_), .B2(new_n1400_), .ZN(new_n1404_));
  INV_X1    g1212(.A(KEYINPUT52), .ZN(new_n1405_));
  OAI21_X1  g1213(.A(new_n1405_), .B1(new_n1219_), .B2(new_n1220_), .ZN(new_n1406_));
  NAND3_X1  g1214(.A1(new_n1207_), .A2(new_n1213_), .A3(KEYINPUT52), .ZN(new_n1407_));
  AND3_X1   g1215(.A1(new_n1406_), .A2(new_n1218_), .A3(new_n1407_), .ZN(new_n1408_));
  AOI21_X1  g1216(.A(new_n1071_), .B1(new_n1221_), .B2(new_n1222_), .ZN(new_n1409_));
  OAI22_X1  g1217(.A1(new_n1402_), .A2(new_n1404_), .B1(new_n1408_), .B2(new_n1409_), .ZN(new_n1410_));
  INV_X1    g1218(.A(new_n1403_), .ZN(new_n1411_));
  NOR3_X1   g1219(.A1(new_n1392_), .A2(new_n1393_), .A3(new_n1249_), .ZN(new_n1412_));
  AOI21_X1  g1220(.A(new_n1398_), .B1(new_n1397_), .B2(new_n1399_), .ZN(new_n1413_));
  OAI21_X1  g1221(.A(new_n1411_), .B1(new_n1412_), .B2(new_n1413_), .ZN(new_n1414_));
  NAND3_X1  g1222(.A1(new_n1406_), .A2(new_n1218_), .A3(new_n1407_), .ZN(new_n1415_));
  NAND3_X1  g1223(.A1(new_n1394_), .A2(new_n1400_), .A3(new_n1403_), .ZN(new_n1416_));
  NAND4_X1  g1224(.A1(new_n1414_), .A2(new_n1216_), .A3(new_n1415_), .A4(new_n1416_), .ZN(new_n1417_));
  NAND2_X1  g1225(.A1(new_n1410_), .A2(new_n1417_), .ZN(new_n1418_));
  INV_X1    g1226(.A(G477gat), .ZN(new_n1419_));
  NOR2_X1   g1227(.A1(new_n205_), .A2(new_n1419_), .ZN(new_n1420_));
  NAND2_X1  g1228(.A1(new_n1418_), .A2(new_n1420_), .ZN(new_n1421_));
  INV_X1    g1229(.A(new_n1420_), .ZN(new_n1422_));
  NAND3_X1  g1230(.A1(new_n1410_), .A2(new_n1422_), .A3(new_n1417_), .ZN(new_n1423_));
  NAND2_X1  g1231(.A1(new_n1421_), .A2(new_n1423_), .ZN(new_n1424_));
  NAND2_X1  g1232(.A1(new_n1248_), .A2(new_n1424_), .ZN(new_n1425_));
  INV_X1    g1233(.A(G494gat), .ZN(new_n1426_));
  NOR2_X1   g1234(.A1(new_n196_), .A2(new_n1426_), .ZN(new_n1427_));
  INV_X1    g1235(.A(new_n1427_), .ZN(new_n1428_));
  NAND3_X1  g1236(.A1(new_n1247_), .A2(new_n1423_), .A3(new_n1421_), .ZN(new_n1429_));
  NAND3_X1  g1237(.A1(new_n1425_), .A2(new_n1428_), .A3(new_n1429_), .ZN(new_n1430_));
  INV_X1    g1238(.A(new_n1430_), .ZN(new_n1431_));
  AOI21_X1  g1239(.A(new_n1428_), .B1(new_n1425_), .B2(new_n1429_), .ZN(new_n1432_));
  NOR2_X1   g1240(.A1(new_n1431_), .A2(new_n1432_), .ZN(new_n1433_));
  NAND3_X1  g1241(.A1(new_n1242_), .A2(new_n1433_), .A3(new_n1236_), .ZN(new_n1434_));
  NAND3_X1  g1242(.A1(new_n1236_), .A2(G1gat), .A3(G494gat), .ZN(new_n1435_));
  NAND2_X1  g1243(.A1(new_n1435_), .A2(new_n1234_), .ZN(new_n1436_));
  OAI21_X1  g1244(.A(new_n1434_), .B1(new_n1433_), .B2(new_n1436_), .ZN(new_n1437_));
  INV_X1    g1245(.A(G511gat), .ZN(new_n1438_));
  NOR2_X1   g1246(.A1(new_n193_), .A2(new_n1438_), .ZN(new_n1439_));
  INV_X1    g1247(.A(new_n1439_), .ZN(new_n1440_));
  XNOR2_X1  g1248(.A(new_n1437_), .B(new_n1440_), .ZN(G5971gat));
  NOR3_X1   g1249(.A1(new_n1436_), .A2(new_n1431_), .A3(new_n1432_), .ZN(new_n1442_));
  AOI21_X1  g1250(.A(new_n1442_), .B1(new_n1437_), .B2(new_n1440_), .ZN(new_n1443_));
  NOR2_X1   g1251(.A1(new_n205_), .A2(new_n1426_), .ZN(new_n1444_));
  AND3_X1   g1252(.A1(new_n1394_), .A2(new_n1400_), .A3(new_n1403_), .ZN(new_n1445_));
  OAI22_X1  g1253(.A1(new_n1445_), .A2(new_n1404_), .B1(new_n1408_), .B2(new_n1409_), .ZN(new_n1446_));
  INV_X1    g1254(.A(KEYINPUT63), .ZN(new_n1447_));
  NAND2_X1  g1255(.A1(new_n1446_), .A2(new_n1447_), .ZN(new_n1448_));
  OAI221_X1 g1256(.A(KEYINPUT63), .B1(new_n1408_), .B2(new_n1409_), .C1(new_n1445_), .C2(new_n1404_), .ZN(new_n1449_));
  AOI22_X1  g1257(.A1(new_n1423_), .A2(KEYINPUT62), .B1(new_n1448_), .B2(new_n1449_), .ZN(new_n1450_));
  INV_X1    g1258(.A(new_n1401_), .ZN(new_n1451_));
  OAI21_X1  g1259(.A(new_n1394_), .B1(new_n1412_), .B2(new_n1451_), .ZN(new_n1452_));
  NAND2_X1  g1260(.A1(new_n1376_), .A2(new_n1378_), .ZN(new_n1453_));
  INV_X1    g1261(.A(new_n1377_), .ZN(new_n1454_));
  NAND2_X1  g1262(.A1(new_n1453_), .A2(new_n1454_), .ZN(new_n1455_));
  NAND3_X1  g1263(.A1(new_n1371_), .A2(new_n1373_), .A3(new_n1375_), .ZN(new_n1456_));
  NAND2_X1  g1264(.A1(new_n1330_), .A2(new_n1333_), .ZN(new_n1457_));
  NAND2_X1  g1265(.A1(new_n1348_), .A2(new_n1457_), .ZN(new_n1458_));
  AOI21_X1  g1266(.A(new_n1261_), .B1(new_n1311_), .B2(new_n1313_), .ZN(new_n1459_));
  OR2_X1    g1267(.A1(new_n1317_), .A2(new_n1459_), .ZN(new_n1460_));
  NOR2_X1   g1268(.A1(new_n944_), .A2(new_n232_), .ZN(new_n1461_));
  NAND2_X1  g1269(.A1(G222gat), .A2(G307gat), .ZN(new_n1462_));
  INV_X1    g1270(.A(new_n1462_), .ZN(new_n1463_));
  NAND2_X1  g1271(.A1(G256gat), .A2(G273gat), .ZN(new_n1464_));
  INV_X1    g1272(.A(new_n1464_), .ZN(new_n1465_));
  NAND3_X1  g1273(.A1(new_n1465_), .A2(new_n1108_), .A3(new_n1268_), .ZN(new_n1466_));
  NAND2_X1  g1274(.A1(G239gat), .A2(G290gat), .ZN(new_n1467_));
  NAND2_X1  g1275(.A1(new_n1467_), .A2(new_n1464_), .ZN(new_n1468_));
  NAND2_X1  g1276(.A1(new_n1466_), .A2(new_n1468_), .ZN(new_n1469_));
  NOR2_X1   g1277(.A1(new_n1465_), .A2(new_n1265_), .ZN(new_n1470_));
  OAI21_X1  g1278(.A(new_n1463_), .B1(new_n1469_), .B2(new_n1470_), .ZN(new_n1471_));
  NAND2_X1  g1279(.A1(new_n1284_), .A2(new_n1464_), .ZN(new_n1472_));
  NAND4_X1  g1280(.A1(new_n1472_), .A2(new_n1466_), .A3(new_n1468_), .A4(new_n1462_), .ZN(new_n1473_));
  NAND2_X1  g1281(.A1(new_n1471_), .A2(new_n1473_), .ZN(new_n1474_));
  INV_X1    g1282(.A(new_n1474_), .ZN(new_n1475_));
  INV_X1    g1283(.A(KEYINPUT65), .ZN(new_n1476_));
  NAND4_X1  g1284(.A1(new_n1286_), .A2(new_n1476_), .A3(new_n1290_), .A4(new_n1287_), .ZN(new_n1477_));
  AND2_X1   g1285(.A1(new_n1477_), .A2(new_n1277_), .ZN(new_n1478_));
  NAND3_X1  g1286(.A1(new_n1286_), .A2(new_n1290_), .A3(new_n1287_), .ZN(new_n1479_));
  NAND2_X1  g1287(.A1(new_n1479_), .A2(KEYINPUT65), .ZN(new_n1480_));
  AOI21_X1  g1288(.A(new_n1475_), .B1(new_n1478_), .B2(new_n1480_), .ZN(new_n1481_));
  INV_X1    g1289(.A(KEYINPUT64), .ZN(new_n1482_));
  AOI21_X1  g1290(.A(new_n1482_), .B1(new_n1471_), .B2(new_n1473_), .ZN(new_n1483_));
  OAI21_X1  g1291(.A(new_n1266_), .B1(new_n1283_), .B2(new_n1290_), .ZN(new_n1484_));
  NOR2_X1   g1292(.A1(new_n1469_), .A2(new_n1470_), .ZN(new_n1485_));
  NAND2_X1  g1293(.A1(new_n1462_), .A2(new_n1482_), .ZN(new_n1486_));
  OAI21_X1  g1294(.A(new_n1484_), .B1(new_n1485_), .B2(new_n1486_), .ZN(new_n1487_));
  NOR2_X1   g1295(.A1(new_n1483_), .A2(new_n1487_), .ZN(new_n1488_));
  OAI21_X1  g1296(.A(new_n1461_), .B1(new_n1481_), .B2(new_n1488_), .ZN(new_n1489_));
  NAND3_X1  g1297(.A1(new_n1480_), .A2(new_n1277_), .A3(new_n1477_), .ZN(new_n1490_));
  NAND2_X1  g1298(.A1(new_n1490_), .A2(new_n1474_), .ZN(new_n1491_));
  INV_X1    g1299(.A(new_n1461_), .ZN(new_n1492_));
  INV_X1    g1300(.A(new_n1488_), .ZN(new_n1493_));
  NAND3_X1  g1301(.A1(new_n1491_), .A2(new_n1492_), .A3(new_n1493_), .ZN(new_n1494_));
  NAND2_X1  g1302(.A1(new_n1489_), .A2(new_n1494_), .ZN(new_n1495_));
  NAND3_X1  g1303(.A1(new_n1293_), .A2(new_n1274_), .A3(new_n1278_), .ZN(new_n1496_));
  AOI22_X1  g1304(.A1(new_n1263_), .A2(new_n1496_), .B1(new_n1295_), .B2(new_n1299_), .ZN(new_n1497_));
  NAND2_X1  g1305(.A1(new_n1495_), .A2(new_n1497_), .ZN(new_n1498_));
  OAI21_X1  g1306(.A(KEYINPUT66), .B1(new_n1481_), .B2(new_n1488_), .ZN(new_n1499_));
  INV_X1    g1307(.A(KEYINPUT66), .ZN(new_n1500_));
  NAND3_X1  g1308(.A1(new_n1491_), .A2(new_n1500_), .A3(new_n1493_), .ZN(new_n1501_));
  AOI21_X1  g1309(.A(new_n1492_), .B1(new_n1499_), .B2(new_n1501_), .ZN(new_n1502_));
  INV_X1    g1310(.A(new_n1497_), .ZN(new_n1503_));
  NAND2_X1  g1311(.A1(new_n1503_), .A2(new_n1494_), .ZN(new_n1504_));
  OAI21_X1  g1312(.A(new_n1498_), .B1(new_n1502_), .B2(new_n1504_), .ZN(new_n1505_));
  NOR2_X1   g1313(.A1(new_n1093_), .A2(new_n258_), .ZN(new_n1506_));
  INV_X1    g1314(.A(new_n1506_), .ZN(new_n1507_));
  NAND2_X1  g1315(.A1(new_n1505_), .A2(new_n1507_), .ZN(new_n1508_));
  NAND2_X1  g1316(.A1(new_n1321_), .A2(new_n1303_), .ZN(new_n1509_));
  NAND2_X1  g1317(.A1(new_n1325_), .A2(new_n1509_), .ZN(new_n1510_));
  OAI211_X1 g1318(.A(new_n1498_), .B(new_n1506_), .C1(new_n1502_), .C2(new_n1504_), .ZN(new_n1511_));
  AND3_X1   g1319(.A1(new_n1508_), .A2(new_n1510_), .A3(new_n1511_), .ZN(new_n1512_));
  AOI21_X1  g1320(.A(new_n1510_), .B1(new_n1508_), .B2(new_n1511_), .ZN(new_n1513_));
  NOR2_X1   g1321(.A1(new_n300_), .A2(new_n799_), .ZN(new_n1514_));
  NOR3_X1   g1322(.A1(new_n1512_), .A2(new_n1513_), .A3(new_n1514_), .ZN(new_n1515_));
  INV_X1    g1323(.A(new_n1514_), .ZN(new_n1516_));
  INV_X1    g1324(.A(new_n1510_), .ZN(new_n1517_));
  INV_X1    g1325(.A(new_n1511_), .ZN(new_n1518_));
  AOI21_X1  g1326(.A(new_n1500_), .B1(new_n1491_), .B2(new_n1493_), .ZN(new_n1519_));
  AOI211_X1 g1327(.A(KEYINPUT66), .B(new_n1488_), .C1(new_n1490_), .C2(new_n1474_), .ZN(new_n1520_));
  OAI21_X1  g1328(.A(new_n1461_), .B1(new_n1519_), .B2(new_n1520_), .ZN(new_n1521_));
  NOR2_X1   g1329(.A1(new_n1481_), .A2(new_n1488_), .ZN(new_n1522_));
  AOI21_X1  g1330(.A(new_n1497_), .B1(new_n1522_), .B2(new_n1492_), .ZN(new_n1523_));
  NAND2_X1  g1331(.A1(new_n1521_), .A2(new_n1523_), .ZN(new_n1524_));
  AOI21_X1  g1332(.A(new_n1506_), .B1(new_n1524_), .B2(new_n1498_), .ZN(new_n1525_));
  OAI21_X1  g1333(.A(new_n1517_), .B1(new_n1518_), .B2(new_n1525_), .ZN(new_n1526_));
  NAND3_X1  g1334(.A1(new_n1508_), .A2(new_n1510_), .A3(new_n1511_), .ZN(new_n1527_));
  AOI21_X1  g1335(.A(new_n1516_), .B1(new_n1526_), .B2(new_n1527_), .ZN(new_n1528_));
  OAI21_X1  g1336(.A(new_n1460_), .B1(new_n1515_), .B2(new_n1528_), .ZN(new_n1529_));
  NOR2_X1   g1337(.A1(new_n960_), .A2(new_n355_), .ZN(new_n1530_));
  INV_X1    g1338(.A(new_n1530_), .ZN(new_n1531_));
  OAI21_X1  g1339(.A(new_n1514_), .B1(new_n1512_), .B2(new_n1513_), .ZN(new_n1532_));
  NOR2_X1   g1340(.A1(new_n1317_), .A2(new_n1459_), .ZN(new_n1533_));
  NAND3_X1  g1341(.A1(new_n1526_), .A2(new_n1516_), .A3(new_n1527_), .ZN(new_n1534_));
  NAND3_X1  g1342(.A1(new_n1532_), .A2(new_n1533_), .A3(new_n1534_), .ZN(new_n1535_));
  AND3_X1   g1343(.A1(new_n1529_), .A2(new_n1531_), .A3(new_n1535_), .ZN(new_n1536_));
  AOI21_X1  g1344(.A(new_n1531_), .B1(new_n1529_), .B2(new_n1535_), .ZN(new_n1537_));
  NOR2_X1   g1345(.A1(new_n1536_), .A2(new_n1537_), .ZN(new_n1538_));
  NAND2_X1  g1346(.A1(new_n1458_), .A2(new_n1538_), .ZN(new_n1539_));
  AND3_X1   g1347(.A1(new_n1532_), .A2(new_n1534_), .A3(new_n1533_), .ZN(new_n1540_));
  AOI21_X1  g1348(.A(new_n1533_), .B1(new_n1532_), .B2(new_n1534_), .ZN(new_n1541_));
  OAI21_X1  g1349(.A(new_n1530_), .B1(new_n1540_), .B2(new_n1541_), .ZN(new_n1542_));
  NAND3_X1  g1350(.A1(new_n1529_), .A2(new_n1531_), .A3(new_n1535_), .ZN(new_n1543_));
  NAND2_X1  g1351(.A1(new_n1542_), .A2(new_n1543_), .ZN(new_n1544_));
  NAND3_X1  g1352(.A1(new_n1544_), .A2(new_n1348_), .A3(new_n1457_), .ZN(new_n1545_));
  NAND2_X1  g1353(.A1(new_n1539_), .A2(new_n1545_), .ZN(new_n1546_));
  NOR2_X1   g1354(.A1(new_n651_), .A2(new_n601_), .ZN(new_n1547_));
  NAND2_X1  g1355(.A1(new_n1546_), .A2(new_n1547_), .ZN(new_n1548_));
  INV_X1    g1356(.A(new_n1547_), .ZN(new_n1549_));
  NAND3_X1  g1357(.A1(new_n1539_), .A2(new_n1549_), .A3(new_n1545_), .ZN(new_n1550_));
  AOI21_X1  g1358(.A(new_n1351_), .B1(new_n1341_), .B2(new_n1350_), .ZN(new_n1551_));
  NOR3_X1   g1359(.A1(new_n1339_), .A2(new_n1340_), .A3(new_n1361_), .ZN(new_n1552_));
  OAI211_X1 g1360(.A(new_n1548_), .B(new_n1550_), .C1(new_n1551_), .C2(new_n1552_), .ZN(new_n1553_));
  OAI21_X1  g1361(.A(new_n1352_), .B1(new_n1360_), .B2(new_n1362_), .ZN(new_n1554_));
  INV_X1    g1362(.A(new_n1552_), .ZN(new_n1555_));
  AND3_X1   g1363(.A1(new_n1539_), .A2(new_n1549_), .A3(new_n1545_), .ZN(new_n1556_));
  AOI21_X1  g1364(.A(new_n1549_), .B1(new_n1539_), .B2(new_n1545_), .ZN(new_n1557_));
  OAI211_X1 g1365(.A(new_n1554_), .B(new_n1555_), .C1(new_n1556_), .C2(new_n1557_), .ZN(new_n1558_));
  NAND2_X1  g1366(.A1(new_n1553_), .A2(new_n1558_), .ZN(new_n1559_));
  NOR2_X1   g1367(.A1(new_n532_), .A2(new_n613_), .ZN(new_n1560_));
  NAND2_X1  g1368(.A1(new_n1559_), .A2(new_n1560_), .ZN(new_n1561_));
  OAI211_X1 g1369(.A(new_n1553_), .B(new_n1558_), .C1(new_n532_), .C2(new_n613_), .ZN(new_n1562_));
  NAND2_X1  g1370(.A1(new_n1561_), .A2(new_n1562_), .ZN(new_n1563_));
  NAND2_X1  g1371(.A1(new_n1363_), .A2(KEYINPUT59), .ZN(new_n1564_));
  NAND2_X1  g1372(.A1(new_n1354_), .A2(new_n1355_), .ZN(new_n1565_));
  NAND3_X1  g1373(.A1(new_n1564_), .A2(new_n1565_), .A3(new_n1353_), .ZN(new_n1566_));
  NAND2_X1  g1374(.A1(new_n1566_), .A2(new_n1253_), .ZN(new_n1567_));
  AOI21_X1  g1375(.A(new_n1366_), .B1(new_n1358_), .B2(new_n1364_), .ZN(new_n1568_));
  INV_X1    g1376(.A(KEYINPUT67), .ZN(new_n1569_));
  OAI21_X1  g1377(.A(new_n1567_), .B1(new_n1568_), .B2(new_n1569_), .ZN(new_n1570_));
  INV_X1    g1378(.A(new_n1364_), .ZN(new_n1571_));
  AOI21_X1  g1379(.A(new_n1571_), .B1(new_n1566_), .B2(new_n1254_), .ZN(new_n1572_));
  NOR3_X1   g1380(.A1(new_n1572_), .A2(KEYINPUT67), .A3(new_n1366_), .ZN(new_n1573_));
  OAI21_X1  g1381(.A(new_n1563_), .B1(new_n1570_), .B2(new_n1573_), .ZN(new_n1574_));
  NAND3_X1  g1382(.A1(new_n1561_), .A2(new_n1562_), .A3(new_n1567_), .ZN(new_n1575_));
  NOR2_X1   g1383(.A1(new_n1575_), .A2(new_n1568_), .ZN(new_n1576_));
  INV_X1    g1384(.A(new_n1576_), .ZN(new_n1577_));
  NOR2_X1   g1385(.A1(new_n452_), .A2(new_n624_), .ZN(new_n1578_));
  AND3_X1   g1386(.A1(new_n1574_), .A2(new_n1577_), .A3(new_n1578_), .ZN(new_n1579_));
  AOI21_X1  g1387(.A(new_n1578_), .B1(new_n1574_), .B2(new_n1577_), .ZN(new_n1580_));
  OAI211_X1 g1388(.A(new_n1455_), .B(new_n1456_), .C1(new_n1579_), .C2(new_n1580_), .ZN(new_n1581_));
  INV_X1    g1389(.A(new_n1578_), .ZN(new_n1582_));
  INV_X1    g1390(.A(new_n1563_), .ZN(new_n1583_));
  INV_X1    g1391(.A(new_n1567_), .ZN(new_n1584_));
  NAND2_X1  g1392(.A1(new_n1365_), .A2(new_n1369_), .ZN(new_n1585_));
  AOI21_X1  g1393(.A(new_n1584_), .B1(new_n1585_), .B2(KEYINPUT67), .ZN(new_n1586_));
  NAND2_X1  g1394(.A1(new_n1568_), .A2(new_n1569_), .ZN(new_n1587_));
  AOI21_X1  g1395(.A(new_n1583_), .B1(new_n1586_), .B2(new_n1587_), .ZN(new_n1588_));
  OAI21_X1  g1396(.A(new_n1582_), .B1(new_n1588_), .B2(new_n1576_), .ZN(new_n1589_));
  OAI21_X1  g1397(.A(KEYINPUT67), .B1(new_n1572_), .B2(new_n1366_), .ZN(new_n1590_));
  NAND3_X1  g1398(.A1(new_n1590_), .A2(new_n1587_), .A3(new_n1567_), .ZN(new_n1591_));
  AOI21_X1  g1399(.A(new_n1576_), .B1(new_n1591_), .B2(new_n1563_), .ZN(new_n1592_));
  NAND2_X1  g1400(.A1(new_n1592_), .A2(new_n1578_), .ZN(new_n1593_));
  INV_X1    g1401(.A(new_n1456_), .ZN(new_n1594_));
  OAI211_X1 g1402(.A(new_n1589_), .B(new_n1593_), .C1(new_n1380_), .C2(new_n1594_), .ZN(new_n1595_));
  NOR2_X1   g1403(.A1(new_n310_), .A2(new_n768_), .ZN(new_n1596_));
  NAND3_X1  g1404(.A1(new_n1581_), .A2(new_n1595_), .A3(new_n1596_), .ZN(new_n1597_));
  NAND2_X1  g1405(.A1(new_n1597_), .A2(KEYINPUT68), .ZN(new_n1598_));
  OAI21_X1  g1406(.A(new_n1387_), .B1(new_n1395_), .B2(new_n1388_), .ZN(new_n1599_));
  INV_X1    g1407(.A(new_n1597_), .ZN(new_n1600_));
  AOI21_X1  g1408(.A(new_n1596_), .B1(new_n1581_), .B2(new_n1595_), .ZN(new_n1601_));
  OAI211_X1 g1409(.A(new_n1598_), .B(new_n1599_), .C1(new_n1600_), .C2(new_n1601_), .ZN(new_n1602_));
  NOR2_X1   g1410(.A1(new_n241_), .A2(new_n918_), .ZN(new_n1603_));
  INV_X1    g1411(.A(new_n1603_), .ZN(new_n1604_));
  NAND2_X1  g1412(.A1(new_n1581_), .A2(new_n1595_), .ZN(new_n1605_));
  INV_X1    g1413(.A(new_n1596_), .ZN(new_n1606_));
  NAND2_X1  g1414(.A1(new_n1605_), .A2(new_n1606_), .ZN(new_n1607_));
  AOI21_X1  g1415(.A(new_n1396_), .B1(new_n1389_), .B2(new_n1391_), .ZN(new_n1608_));
  OAI211_X1 g1416(.A(new_n1597_), .B(new_n1607_), .C1(new_n1608_), .C2(KEYINPUT68), .ZN(new_n1609_));
  AND3_X1   g1417(.A1(new_n1602_), .A2(new_n1604_), .A3(new_n1609_), .ZN(new_n1610_));
  AOI21_X1  g1418(.A(new_n1604_), .B1(new_n1602_), .B2(new_n1609_), .ZN(new_n1611_));
  OAI21_X1  g1419(.A(new_n1452_), .B1(new_n1610_), .B2(new_n1611_), .ZN(new_n1612_));
  NAND2_X1  g1420(.A1(new_n1602_), .A2(new_n1609_), .ZN(new_n1613_));
  NAND2_X1  g1421(.A1(new_n1613_), .A2(new_n1603_), .ZN(new_n1614_));
  NAND3_X1  g1422(.A1(new_n1602_), .A2(new_n1604_), .A3(new_n1609_), .ZN(new_n1615_));
  AOI21_X1  g1423(.A(new_n1413_), .B1(new_n1400_), .B2(new_n1403_), .ZN(new_n1616_));
  NAND3_X1  g1424(.A1(new_n1614_), .A2(new_n1615_), .A3(new_n1616_), .ZN(new_n1617_));
  NOR2_X1   g1425(.A1(new_n215_), .A2(new_n1419_), .ZN(new_n1618_));
  INV_X1    g1426(.A(new_n1618_), .ZN(new_n1619_));
  NAND3_X1  g1427(.A1(new_n1612_), .A2(new_n1617_), .A3(new_n1619_), .ZN(new_n1620_));
  NAND2_X1  g1428(.A1(new_n1612_), .A2(new_n1617_), .ZN(new_n1621_));
  NAND2_X1  g1429(.A1(new_n1621_), .A2(new_n1618_), .ZN(new_n1622_));
  INV_X1    g1430(.A(KEYINPUT62), .ZN(new_n1623_));
  NAND4_X1  g1431(.A1(new_n1410_), .A2(new_n1417_), .A3(new_n1623_), .A4(new_n1422_), .ZN(new_n1624_));
  NAND4_X1  g1432(.A1(new_n1450_), .A2(new_n1620_), .A3(new_n1622_), .A4(new_n1624_), .ZN(new_n1625_));
  NAND2_X1  g1433(.A1(new_n1423_), .A2(new_n1446_), .ZN(new_n1626_));
  AND3_X1   g1434(.A1(new_n1612_), .A2(new_n1617_), .A3(new_n1619_), .ZN(new_n1627_));
  AOI21_X1  g1435(.A(new_n1619_), .B1(new_n1612_), .B2(new_n1617_), .ZN(new_n1628_));
  OAI21_X1  g1436(.A(new_n1626_), .B1(new_n1627_), .B2(new_n1628_), .ZN(new_n1629_));
  AOI21_X1  g1437(.A(new_n1444_), .B1(new_n1625_), .B2(new_n1629_), .ZN(new_n1630_));
  NAND2_X1  g1438(.A1(new_n1423_), .A2(KEYINPUT62), .ZN(new_n1631_));
  NAND2_X1  g1439(.A1(new_n1448_), .A2(new_n1449_), .ZN(new_n1632_));
  NAND3_X1  g1440(.A1(new_n1631_), .A2(new_n1632_), .A3(new_n1624_), .ZN(new_n1633_));
  NAND2_X1  g1441(.A1(new_n1622_), .A2(new_n1620_), .ZN(new_n1634_));
  OAI211_X1 g1442(.A(new_n1629_), .B(new_n1444_), .C1(new_n1633_), .C2(new_n1634_), .ZN(new_n1635_));
  INV_X1    g1443(.A(new_n1635_), .ZN(new_n1636_));
  OAI211_X1 g1444(.A(new_n1429_), .B(new_n1430_), .C1(new_n1630_), .C2(new_n1636_), .ZN(new_n1637_));
  OAI21_X1  g1445(.A(new_n1629_), .B1(new_n1633_), .B2(new_n1634_), .ZN(new_n1638_));
  INV_X1    g1446(.A(new_n1444_), .ZN(new_n1639_));
  NAND2_X1  g1447(.A1(new_n1638_), .A2(new_n1639_), .ZN(new_n1640_));
  AOI21_X1  g1448(.A(new_n1247_), .B1(new_n1423_), .B2(new_n1421_), .ZN(new_n1641_));
  OAI21_X1  g1449(.A(new_n1429_), .B1(new_n1641_), .B2(new_n1427_), .ZN(new_n1642_));
  NAND3_X1  g1450(.A1(new_n1640_), .A2(new_n1642_), .A3(new_n1635_), .ZN(new_n1643_));
  NAND2_X1  g1451(.A1(new_n1637_), .A2(new_n1643_), .ZN(new_n1644_));
  NOR2_X1   g1452(.A1(new_n196_), .A2(new_n1438_), .ZN(new_n1645_));
  NAND2_X1  g1453(.A1(new_n1644_), .A2(new_n1645_), .ZN(new_n1646_));
  INV_X1    g1454(.A(new_n1645_), .ZN(new_n1647_));
  NAND3_X1  g1455(.A1(new_n1637_), .A2(new_n1647_), .A3(new_n1643_), .ZN(new_n1648_));
  NAND2_X1  g1456(.A1(new_n1646_), .A2(new_n1648_), .ZN(new_n1649_));
  NOR2_X1   g1457(.A1(new_n1443_), .A2(new_n1649_), .ZN(new_n1650_));
  INV_X1    g1458(.A(new_n1650_), .ZN(new_n1651_));
  NAND2_X1  g1459(.A1(new_n1443_), .A2(new_n1649_), .ZN(new_n1652_));
  NAND2_X1  g1460(.A1(new_n1651_), .A2(new_n1652_), .ZN(new_n1653_));
  INV_X1    g1461(.A(G528gat), .ZN(new_n1654_));
  NOR2_X1   g1462(.A1(new_n193_), .A2(new_n1654_), .ZN(new_n1655_));
  XNOR2_X1  g1463(.A(new_n1653_), .B(new_n1655_), .ZN(G6123gat));
  INV_X1    g1464(.A(new_n1655_), .ZN(new_n1657_));
  AOI21_X1  g1465(.A(new_n1650_), .B1(new_n1657_), .B2(new_n1652_), .ZN(new_n1658_));
  NAND3_X1  g1466(.A1(new_n1622_), .A2(new_n1626_), .A3(new_n1620_), .ZN(new_n1659_));
  NAND2_X1  g1467(.A1(new_n1640_), .A2(new_n1659_), .ZN(new_n1660_));
  OR3_X1    g1468(.A1(new_n1610_), .A2(new_n1611_), .A3(new_n1452_), .ZN(new_n1661_));
  OAI21_X1  g1469(.A(new_n1599_), .B1(new_n1600_), .B2(new_n1601_), .ZN(new_n1662_));
  NAND2_X1  g1470(.A1(new_n1615_), .A2(new_n1662_), .ZN(new_n1663_));
  NAND2_X1  g1471(.A1(new_n1595_), .A2(new_n1596_), .ZN(new_n1664_));
  NAND2_X1  g1472(.A1(new_n1664_), .A2(new_n1581_), .ZN(new_n1665_));
  NOR2_X1   g1473(.A1(new_n532_), .A2(new_n624_), .ZN(new_n1666_));
  NOR2_X1   g1474(.A1(new_n1458_), .A2(new_n1538_), .ZN(new_n1667_));
  OAI21_X1  g1475(.A(new_n1539_), .B1(new_n1667_), .B2(new_n1547_), .ZN(new_n1668_));
  AOI21_X1  g1476(.A(new_n1540_), .B1(new_n1531_), .B2(new_n1529_), .ZN(new_n1669_));
  AOI21_X1  g1477(.A(new_n1512_), .B1(new_n1516_), .B2(new_n1526_), .ZN(new_n1670_));
  AOI22_X1  g1478(.A1(new_n1505_), .A2(new_n1507_), .B1(new_n1503_), .B2(new_n1495_), .ZN(new_n1671_));
  OR2_X1    g1479(.A1(new_n1469_), .A2(KEYINPUT70), .ZN(new_n1672_));
  NAND2_X1  g1480(.A1(new_n1469_), .A2(KEYINPUT70), .ZN(new_n1673_));
  NAND3_X1  g1481(.A1(new_n1672_), .A2(new_n1473_), .A3(new_n1673_), .ZN(new_n1674_));
  NAND3_X1  g1482(.A1(new_n1270_), .A2(G256gat), .A3(G290gat), .ZN(new_n1675_));
  INV_X1    g1483(.A(G239gat), .ZN(new_n1676_));
  NOR2_X1   g1484(.A1(new_n1676_), .A2(new_n211_), .ZN(new_n1677_));
  XNOR2_X1  g1485(.A(new_n1675_), .B(new_n1677_), .ZN(new_n1678_));
  INV_X1    g1486(.A(new_n1678_), .ZN(new_n1679_));
  NAND2_X1  g1487(.A1(new_n1674_), .A2(new_n1679_), .ZN(new_n1680_));
  INV_X1    g1488(.A(G222gat), .ZN(new_n1681_));
  NOR2_X1   g1489(.A1(new_n1681_), .A2(new_n232_), .ZN(new_n1682_));
  INV_X1    g1490(.A(new_n1682_), .ZN(new_n1683_));
  OAI211_X1 g1491(.A(new_n1468_), .B(new_n1466_), .C1(new_n1470_), .C2(new_n1463_), .ZN(new_n1684_));
  OAI211_X1 g1492(.A(new_n1680_), .B(new_n1683_), .C1(new_n1679_), .C2(new_n1684_), .ZN(new_n1685_));
  NOR2_X1   g1493(.A1(new_n1684_), .A2(new_n1678_), .ZN(new_n1686_));
  AOI21_X1  g1494(.A(new_n1686_), .B1(new_n1674_), .B2(new_n1678_), .ZN(new_n1687_));
  NAND2_X1  g1495(.A1(new_n1687_), .A2(new_n1682_), .ZN(new_n1688_));
  NAND2_X1  g1496(.A1(new_n1685_), .A2(new_n1688_), .ZN(new_n1689_));
  OAI21_X1  g1497(.A(new_n1492_), .B1(new_n1519_), .B2(new_n1520_), .ZN(new_n1690_));
  NOR2_X1   g1498(.A1(new_n1474_), .A2(new_n1484_), .ZN(new_n1691_));
  INV_X1    g1499(.A(new_n1691_), .ZN(new_n1692_));
  AOI21_X1  g1500(.A(new_n1689_), .B1(new_n1690_), .B2(new_n1692_), .ZN(new_n1693_));
  OAI211_X1 g1501(.A(new_n1692_), .B(new_n1689_), .C1(new_n1522_), .C2(new_n1461_), .ZN(new_n1694_));
  INV_X1    g1502(.A(new_n1694_), .ZN(new_n1695_));
  NOR2_X1   g1503(.A1(new_n944_), .A2(new_n258_), .ZN(new_n1696_));
  NOR3_X1   g1504(.A1(new_n1693_), .A2(new_n1695_), .A3(new_n1696_), .ZN(new_n1697_));
  INV_X1    g1505(.A(new_n1696_), .ZN(new_n1698_));
  INV_X1    g1506(.A(new_n1689_), .ZN(new_n1699_));
  AOI21_X1  g1507(.A(new_n1461_), .B1(new_n1499_), .B2(new_n1501_), .ZN(new_n1700_));
  OAI21_X1  g1508(.A(new_n1699_), .B1(new_n1700_), .B2(new_n1691_), .ZN(new_n1701_));
  AOI21_X1  g1509(.A(new_n1698_), .B1(new_n1701_), .B2(new_n1694_), .ZN(new_n1702_));
  OAI21_X1  g1510(.A(new_n1671_), .B1(new_n1697_), .B2(new_n1702_), .ZN(new_n1703_));
  NAND2_X1  g1511(.A1(new_n1495_), .A2(new_n1503_), .ZN(new_n1704_));
  AOI22_X1  g1512(.A1(new_n1521_), .A2(new_n1523_), .B1(new_n1497_), .B2(new_n1495_), .ZN(new_n1705_));
  OAI21_X1  g1513(.A(new_n1704_), .B1(new_n1705_), .B2(new_n1506_), .ZN(new_n1706_));
  OAI21_X1  g1514(.A(new_n1696_), .B1(new_n1693_), .B2(new_n1695_), .ZN(new_n1707_));
  NAND3_X1  g1515(.A1(new_n1701_), .A2(new_n1698_), .A3(new_n1694_), .ZN(new_n1708_));
  NAND3_X1  g1516(.A1(new_n1706_), .A2(new_n1707_), .A3(new_n1708_), .ZN(new_n1709_));
  NOR2_X1   g1517(.A1(new_n300_), .A2(new_n1093_), .ZN(new_n1710_));
  INV_X1    g1518(.A(new_n1710_), .ZN(new_n1711_));
  AND3_X1   g1519(.A1(new_n1703_), .A2(new_n1709_), .A3(new_n1711_), .ZN(new_n1712_));
  AOI21_X1  g1520(.A(new_n1711_), .B1(new_n1703_), .B2(new_n1709_), .ZN(new_n1713_));
  OAI21_X1  g1521(.A(new_n1670_), .B1(new_n1712_), .B2(new_n1713_), .ZN(new_n1714_));
  NAND2_X1  g1522(.A1(new_n1703_), .A2(new_n1709_), .ZN(new_n1715_));
  NAND2_X1  g1523(.A1(new_n1715_), .A2(new_n1710_), .ZN(new_n1716_));
  NAND2_X1  g1524(.A1(new_n1534_), .A2(new_n1527_), .ZN(new_n1717_));
  NAND3_X1  g1525(.A1(new_n1703_), .A2(new_n1709_), .A3(new_n1711_), .ZN(new_n1718_));
  NAND3_X1  g1526(.A1(new_n1716_), .A2(new_n1717_), .A3(new_n1718_), .ZN(new_n1719_));
  NOR2_X1   g1527(.A1(new_n799_), .A2(new_n355_), .ZN(new_n1720_));
  INV_X1    g1528(.A(new_n1720_), .ZN(new_n1721_));
  NAND3_X1  g1529(.A1(new_n1714_), .A2(new_n1719_), .A3(new_n1721_), .ZN(new_n1722_));
  INV_X1    g1530(.A(new_n1722_), .ZN(new_n1723_));
  AOI21_X1  g1531(.A(new_n1721_), .B1(new_n1714_), .B2(new_n1719_), .ZN(new_n1724_));
  OAI21_X1  g1532(.A(new_n1669_), .B1(new_n1723_), .B2(new_n1724_), .ZN(new_n1725_));
  NAND2_X1  g1533(.A1(new_n1714_), .A2(new_n1719_), .ZN(new_n1726_));
  NAND2_X1  g1534(.A1(new_n1726_), .A2(new_n1720_), .ZN(new_n1727_));
  OAI21_X1  g1535(.A(new_n1535_), .B1(new_n1541_), .B2(new_n1530_), .ZN(new_n1728_));
  NAND3_X1  g1536(.A1(new_n1727_), .A2(new_n1728_), .A3(new_n1722_), .ZN(new_n1729_));
  NOR2_X1   g1537(.A1(new_n960_), .A2(new_n601_), .ZN(new_n1730_));
  INV_X1    g1538(.A(new_n1730_), .ZN(new_n1731_));
  NAND3_X1  g1539(.A1(new_n1725_), .A2(new_n1729_), .A3(new_n1731_), .ZN(new_n1732_));
  INV_X1    g1540(.A(new_n1732_), .ZN(new_n1733_));
  AOI21_X1  g1541(.A(new_n1731_), .B1(new_n1725_), .B2(new_n1729_), .ZN(new_n1734_));
  OAI21_X1  g1542(.A(new_n1668_), .B1(new_n1733_), .B2(new_n1734_), .ZN(new_n1735_));
  NOR3_X1   g1543(.A1(new_n1723_), .A2(new_n1724_), .A3(new_n1669_), .ZN(new_n1736_));
  AOI21_X1  g1544(.A(new_n1728_), .B1(new_n1727_), .B2(new_n1722_), .ZN(new_n1737_));
  OAI21_X1  g1545(.A(new_n1730_), .B1(new_n1736_), .B2(new_n1737_), .ZN(new_n1738_));
  NAND4_X1  g1546(.A1(new_n1738_), .A2(new_n1550_), .A3(new_n1732_), .A4(new_n1539_), .ZN(new_n1739_));
  NAND2_X1  g1547(.A1(G137gat), .A2(G409gat), .ZN(new_n1740_));
  NAND3_X1  g1548(.A1(new_n1735_), .A2(new_n1739_), .A3(new_n1740_), .ZN(new_n1741_));
  INV_X1    g1549(.A(new_n1741_), .ZN(new_n1742_));
  AOI21_X1  g1550(.A(new_n1740_), .B1(new_n1735_), .B2(new_n1739_), .ZN(new_n1743_));
  OAI211_X1 g1551(.A(new_n1562_), .B(new_n1553_), .C1(new_n1742_), .C2(new_n1743_), .ZN(new_n1744_));
  INV_X1    g1552(.A(new_n1558_), .ZN(new_n1745_));
  OAI21_X1  g1553(.A(new_n1553_), .B1(new_n1745_), .B2(new_n1560_), .ZN(new_n1746_));
  INV_X1    g1554(.A(new_n1743_), .ZN(new_n1747_));
  INV_X1    g1555(.A(KEYINPUT71), .ZN(new_n1748_));
  NAND2_X1  g1556(.A1(new_n1741_), .A2(new_n1748_), .ZN(new_n1749_));
  NAND4_X1  g1557(.A1(new_n1735_), .A2(new_n1739_), .A3(KEYINPUT71), .A4(new_n1740_), .ZN(new_n1750_));
  NAND4_X1  g1558(.A1(new_n1746_), .A2(new_n1747_), .A3(new_n1749_), .A4(new_n1750_), .ZN(new_n1751_));
  INV_X1    g1559(.A(KEYINPUT72), .ZN(new_n1752_));
  OAI21_X1  g1560(.A(new_n1744_), .B1(new_n1751_), .B2(new_n1752_), .ZN(new_n1753_));
  AND2_X1   g1561(.A1(new_n1749_), .A2(new_n1750_), .ZN(new_n1754_));
  AOI21_X1  g1562(.A(new_n1743_), .B1(new_n1562_), .B2(new_n1553_), .ZN(new_n1755_));
  AOI21_X1  g1563(.A(KEYINPUT72), .B1(new_n1754_), .B2(new_n1755_), .ZN(new_n1756_));
  OAI21_X1  g1564(.A(new_n1666_), .B1(new_n1753_), .B2(new_n1756_), .ZN(new_n1757_));
  NAND3_X1  g1565(.A1(new_n1754_), .A2(new_n1755_), .A3(KEYINPUT72), .ZN(new_n1758_));
  NAND2_X1  g1566(.A1(new_n1751_), .A2(new_n1752_), .ZN(new_n1759_));
  INV_X1    g1567(.A(new_n1666_), .ZN(new_n1760_));
  NAND4_X1  g1568(.A1(new_n1758_), .A2(new_n1759_), .A3(new_n1760_), .A4(new_n1744_), .ZN(new_n1761_));
  AND2_X1   g1569(.A1(new_n1757_), .A2(new_n1761_), .ZN(new_n1762_));
  NAND2_X1  g1570(.A1(new_n1574_), .A2(new_n1577_), .ZN(new_n1763_));
  AOI22_X1  g1571(.A1(new_n1763_), .A2(new_n1582_), .B1(new_n1583_), .B2(new_n1591_), .ZN(new_n1764_));
  NAND3_X1  g1572(.A1(new_n1758_), .A2(new_n1759_), .A3(new_n1744_), .ZN(new_n1765_));
  AOI21_X1  g1573(.A(KEYINPUT73), .B1(new_n1765_), .B2(new_n1666_), .ZN(new_n1766_));
  OAI21_X1  g1574(.A(new_n1762_), .B1(new_n1764_), .B2(new_n1766_), .ZN(new_n1767_));
  NOR2_X1   g1575(.A1(new_n452_), .A2(new_n768_), .ZN(new_n1768_));
  INV_X1    g1576(.A(new_n1768_), .ZN(new_n1769_));
  NAND2_X1  g1577(.A1(new_n1591_), .A2(new_n1583_), .ZN(new_n1770_));
  OAI21_X1  g1578(.A(new_n1770_), .B1(new_n1592_), .B2(new_n1578_), .ZN(new_n1771_));
  INV_X1    g1579(.A(KEYINPUT73), .ZN(new_n1772_));
  NAND2_X1  g1580(.A1(new_n1757_), .A2(new_n1772_), .ZN(new_n1773_));
  NAND2_X1  g1581(.A1(new_n1757_), .A2(new_n1761_), .ZN(new_n1774_));
  NAND3_X1  g1582(.A1(new_n1771_), .A2(new_n1773_), .A3(new_n1774_), .ZN(new_n1775_));
  AND3_X1   g1583(.A1(new_n1767_), .A2(new_n1769_), .A3(new_n1775_), .ZN(new_n1776_));
  AOI21_X1  g1584(.A(new_n1769_), .B1(new_n1767_), .B2(new_n1775_), .ZN(new_n1777_));
  OAI21_X1  g1585(.A(new_n1665_), .B1(new_n1776_), .B2(new_n1777_), .ZN(new_n1778_));
  NOR2_X1   g1586(.A1(new_n310_), .A2(new_n918_), .ZN(new_n1779_));
  INV_X1    g1587(.A(new_n1779_), .ZN(new_n1780_));
  NOR2_X1   g1588(.A1(new_n1579_), .A2(new_n1580_), .ZN(new_n1781_));
  NAND2_X1  g1589(.A1(new_n1455_), .A2(new_n1456_), .ZN(new_n1782_));
  AOI21_X1  g1590(.A(new_n1606_), .B1(new_n1781_), .B2(new_n1782_), .ZN(new_n1783_));
  INV_X1    g1591(.A(new_n1581_), .ZN(new_n1784_));
  NOR2_X1   g1592(.A1(new_n1783_), .A2(new_n1784_), .ZN(new_n1785_));
  AND3_X1   g1593(.A1(new_n1771_), .A2(new_n1773_), .A3(new_n1774_), .ZN(new_n1786_));
  AOI21_X1  g1594(.A(new_n1774_), .B1(new_n1771_), .B2(new_n1773_), .ZN(new_n1787_));
  OAI21_X1  g1595(.A(new_n1768_), .B1(new_n1786_), .B2(new_n1787_), .ZN(new_n1788_));
  NAND3_X1  g1596(.A1(new_n1767_), .A2(new_n1769_), .A3(new_n1775_), .ZN(new_n1789_));
  NAND3_X1  g1597(.A1(new_n1785_), .A2(new_n1788_), .A3(new_n1789_), .ZN(new_n1790_));
  NAND3_X1  g1598(.A1(new_n1778_), .A2(new_n1780_), .A3(new_n1790_), .ZN(new_n1791_));
  AOI21_X1  g1599(.A(new_n1780_), .B1(new_n1778_), .B2(new_n1790_), .ZN(new_n1792_));
  INV_X1    g1600(.A(new_n1792_), .ZN(new_n1793_));
  NAND3_X1  g1601(.A1(new_n1663_), .A2(new_n1791_), .A3(new_n1793_), .ZN(new_n1794_));
  NOR2_X1   g1602(.A1(new_n241_), .A2(new_n1419_), .ZN(new_n1795_));
  INV_X1    g1603(.A(new_n1795_), .ZN(new_n1796_));
  AND3_X1   g1604(.A1(new_n1778_), .A2(new_n1780_), .A3(new_n1790_), .ZN(new_n1797_));
  OAI211_X1 g1605(.A(new_n1615_), .B(new_n1662_), .C1(new_n1797_), .C2(new_n1792_), .ZN(new_n1798_));
  AND3_X1   g1606(.A1(new_n1794_), .A2(new_n1796_), .A3(new_n1798_), .ZN(new_n1799_));
  AOI21_X1  g1607(.A(new_n1796_), .B1(new_n1794_), .B2(new_n1798_), .ZN(new_n1800_));
  OAI211_X1 g1608(.A(new_n1620_), .B(new_n1661_), .C1(new_n1799_), .C2(new_n1800_), .ZN(new_n1801_));
  NAND2_X1  g1609(.A1(new_n1620_), .A2(new_n1661_), .ZN(new_n1802_));
  NAND2_X1  g1610(.A1(new_n1794_), .A2(new_n1798_), .ZN(new_n1803_));
  NAND2_X1  g1611(.A1(new_n1803_), .A2(new_n1795_), .ZN(new_n1804_));
  NAND3_X1  g1612(.A1(new_n1794_), .A2(new_n1798_), .A3(new_n1796_), .ZN(new_n1805_));
  NAND3_X1  g1613(.A1(new_n1802_), .A2(new_n1804_), .A3(new_n1805_), .ZN(new_n1806_));
  NAND2_X1  g1614(.A1(new_n1801_), .A2(new_n1806_), .ZN(new_n1807_));
  NOR2_X1   g1615(.A1(new_n215_), .A2(new_n1426_), .ZN(new_n1808_));
  INV_X1    g1616(.A(new_n1808_), .ZN(new_n1809_));
  NAND2_X1  g1617(.A1(new_n1807_), .A2(new_n1809_), .ZN(new_n1810_));
  NAND3_X1  g1618(.A1(new_n1801_), .A2(new_n1806_), .A3(new_n1808_), .ZN(new_n1811_));
  NAND2_X1  g1619(.A1(new_n1810_), .A2(new_n1811_), .ZN(new_n1812_));
  INV_X1    g1620(.A(KEYINPUT74), .ZN(new_n1813_));
  NAND2_X1  g1621(.A1(new_n1811_), .A2(new_n1813_), .ZN(new_n1814_));
  NAND3_X1  g1622(.A1(new_n1660_), .A2(new_n1812_), .A3(new_n1814_), .ZN(new_n1815_));
  INV_X1    g1623(.A(new_n1659_), .ZN(new_n1816_));
  AOI21_X1  g1624(.A(new_n1816_), .B1(new_n1638_), .B2(new_n1639_), .ZN(new_n1817_));
  OAI211_X1 g1625(.A(new_n1811_), .B(new_n1810_), .C1(new_n1817_), .C2(new_n1813_), .ZN(new_n1818_));
  NAND2_X1  g1626(.A1(new_n1815_), .A2(new_n1818_), .ZN(new_n1819_));
  NOR2_X1   g1627(.A1(new_n205_), .A2(new_n1438_), .ZN(new_n1820_));
  NAND2_X1  g1628(.A1(new_n1819_), .A2(new_n1820_), .ZN(new_n1821_));
  OAI21_X1  g1629(.A(KEYINPUT69), .B1(new_n1630_), .B2(new_n1636_), .ZN(new_n1822_));
  INV_X1    g1630(.A(KEYINPUT69), .ZN(new_n1823_));
  NAND3_X1  g1631(.A1(new_n1640_), .A2(new_n1823_), .A3(new_n1635_), .ZN(new_n1824_));
  NAND3_X1  g1632(.A1(new_n1822_), .A2(new_n1642_), .A3(new_n1824_), .ZN(new_n1825_));
  NAND2_X1  g1633(.A1(new_n1648_), .A2(new_n1825_), .ZN(new_n1826_));
  INV_X1    g1634(.A(new_n1820_), .ZN(new_n1827_));
  NAND3_X1  g1635(.A1(new_n1815_), .A2(new_n1818_), .A3(new_n1827_), .ZN(new_n1828_));
  AND3_X1   g1636(.A1(new_n1821_), .A2(new_n1826_), .A3(new_n1828_), .ZN(new_n1829_));
  AOI21_X1  g1637(.A(new_n1826_), .B1(new_n1828_), .B2(new_n1821_), .ZN(new_n1830_));
  NOR2_X1   g1638(.A1(new_n196_), .A2(new_n1654_), .ZN(new_n1831_));
  NOR3_X1   g1639(.A1(new_n1829_), .A2(new_n1830_), .A3(new_n1831_), .ZN(new_n1832_));
  INV_X1    g1640(.A(new_n1831_), .ZN(new_n1833_));
  NAND2_X1  g1641(.A1(new_n1821_), .A2(new_n1828_), .ZN(new_n1834_));
  INV_X1    g1642(.A(new_n1826_), .ZN(new_n1835_));
  NAND2_X1  g1643(.A1(new_n1834_), .A2(new_n1835_), .ZN(new_n1836_));
  NAND3_X1  g1644(.A1(new_n1821_), .A2(new_n1826_), .A3(new_n1828_), .ZN(new_n1837_));
  AOI21_X1  g1645(.A(new_n1833_), .B1(new_n1836_), .B2(new_n1837_), .ZN(new_n1838_));
  OAI21_X1  g1646(.A(new_n1658_), .B1(new_n1832_), .B2(new_n1838_), .ZN(new_n1839_));
  INV_X1    g1647(.A(new_n1839_), .ZN(new_n1840_));
  NOR3_X1   g1648(.A1(new_n1658_), .A2(new_n1832_), .A3(new_n1838_), .ZN(new_n1841_));
  NOR2_X1   g1649(.A1(new_n1840_), .A2(new_n1841_), .ZN(G6150gat));
  AOI21_X1  g1650(.A(new_n1829_), .B1(new_n1836_), .B2(new_n1833_), .ZN(new_n1843_));
  NAND2_X1  g1651(.A1(new_n1660_), .A2(new_n1812_), .ZN(new_n1844_));
  NAND3_X1  g1652(.A1(new_n1801_), .A2(new_n1806_), .A3(new_n1809_), .ZN(new_n1845_));
  NAND2_X1  g1653(.A1(new_n1845_), .A2(KEYINPUT75), .ZN(new_n1846_));
  INV_X1    g1654(.A(new_n1790_), .ZN(new_n1847_));
  AOI21_X1  g1655(.A(new_n1847_), .B1(new_n1780_), .B2(new_n1778_), .ZN(new_n1848_));
  NAND2_X1  g1656(.A1(new_n1747_), .A2(new_n1741_), .ZN(new_n1849_));
  NAND2_X1  g1657(.A1(new_n1849_), .A2(new_n1746_), .ZN(new_n1850_));
  INV_X1    g1658(.A(new_n1850_), .ZN(new_n1851_));
  OAI21_X1  g1659(.A(new_n1760_), .B1(new_n1753_), .B2(new_n1756_), .ZN(new_n1852_));
  AOI21_X1  g1660(.A(new_n1851_), .B1(new_n1852_), .B2(KEYINPUT82), .ZN(new_n1853_));
  INV_X1    g1661(.A(KEYINPUT82), .ZN(new_n1854_));
  NAND3_X1  g1662(.A1(new_n1765_), .A2(new_n1854_), .A3(new_n1760_), .ZN(new_n1855_));
  NAND2_X1  g1663(.A1(new_n1853_), .A2(new_n1855_), .ZN(new_n1856_));
  NOR2_X1   g1664(.A1(new_n651_), .A2(new_n624_), .ZN(new_n1857_));
  INV_X1    g1665(.A(KEYINPUT78), .ZN(new_n1858_));
  OAI211_X1 g1666(.A(new_n1732_), .B(new_n1738_), .C1(new_n1668_), .C2(new_n1858_), .ZN(new_n1859_));
  NAND3_X1  g1667(.A1(new_n1859_), .A2(G137gat), .A3(G409gat), .ZN(new_n1860_));
  NAND2_X1  g1668(.A1(new_n1668_), .A2(KEYINPUT78), .ZN(new_n1861_));
  NAND3_X1  g1669(.A1(new_n1735_), .A2(new_n1739_), .A3(new_n1861_), .ZN(new_n1862_));
  NAND2_X1  g1670(.A1(new_n1860_), .A2(new_n1862_), .ZN(new_n1863_));
  INV_X1    g1671(.A(new_n1863_), .ZN(new_n1864_));
  AOI21_X1  g1672(.A(new_n1736_), .B1(new_n1731_), .B2(new_n1725_), .ZN(new_n1865_));
  NOR2_X1   g1673(.A1(new_n799_), .A2(new_n601_), .ZN(new_n1866_));
  INV_X1    g1674(.A(new_n1866_), .ZN(new_n1867_));
  AOI21_X1  g1675(.A(new_n1706_), .B1(new_n1708_), .B2(new_n1707_), .ZN(new_n1868_));
  OAI21_X1  g1676(.A(new_n1709_), .B1(new_n1868_), .B2(new_n1710_), .ZN(new_n1869_));
  OAI21_X1  g1677(.A(new_n1701_), .B1(new_n1695_), .B2(new_n1696_), .ZN(new_n1870_));
  OAI21_X1  g1678(.A(new_n1683_), .B1(new_n1679_), .B2(new_n1684_), .ZN(new_n1871_));
  INV_X1    g1679(.A(G256gat), .ZN(new_n1872_));
  NAND2_X1  g1680(.A1(new_n1268_), .A2(G273gat), .ZN(new_n1873_));
  AOI21_X1  g1681(.A(new_n1872_), .B1(new_n1873_), .B2(new_n211_), .ZN(new_n1874_));
  NAND2_X1  g1682(.A1(new_n1677_), .A2(G290gat), .ZN(new_n1875_));
  NAND2_X1  g1683(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1876_));
  NAND2_X1  g1684(.A1(G239gat), .A2(G324gat), .ZN(new_n1877_));
  XNOR2_X1  g1685(.A(new_n1876_), .B(new_n1877_), .ZN(new_n1878_));
  AND3_X1   g1686(.A1(new_n1680_), .A2(new_n1871_), .A3(new_n1878_), .ZN(new_n1879_));
  OAI21_X1  g1687(.A(new_n1680_), .B1(new_n1687_), .B2(new_n1682_), .ZN(new_n1880_));
  INV_X1    g1688(.A(new_n1878_), .ZN(new_n1881_));
  AOI21_X1  g1689(.A(new_n1879_), .B1(new_n1880_), .B2(new_n1881_), .ZN(new_n1882_));
  NOR2_X1   g1690(.A1(new_n1681_), .A2(new_n258_), .ZN(new_n1883_));
  AND2_X1   g1691(.A1(new_n1680_), .A2(new_n1871_), .ZN(new_n1884_));
  AOI21_X1  g1692(.A(new_n1883_), .B1(new_n1884_), .B2(new_n1881_), .ZN(new_n1885_));
  NAND2_X1  g1693(.A1(new_n1880_), .A2(new_n1878_), .ZN(new_n1886_));
  AOI22_X1  g1694(.A1(new_n1882_), .A2(new_n1883_), .B1(new_n1885_), .B2(new_n1886_), .ZN(new_n1887_));
  NAND2_X1  g1695(.A1(new_n1870_), .A2(new_n1887_), .ZN(new_n1888_));
  NAND2_X1  g1696(.A1(new_n1690_), .A2(new_n1692_), .ZN(new_n1889_));
  AOI22_X1  g1697(.A1(new_n1889_), .A2(new_n1699_), .B1(new_n1698_), .B2(new_n1694_), .ZN(new_n1890_));
  INV_X1    g1698(.A(new_n1887_), .ZN(new_n1891_));
  NAND2_X1  g1699(.A1(new_n1890_), .A2(new_n1891_), .ZN(new_n1892_));
  NOR2_X1   g1700(.A1(new_n300_), .A2(new_n944_), .ZN(new_n1893_));
  INV_X1    g1701(.A(new_n1893_), .ZN(new_n1894_));
  NAND3_X1  g1702(.A1(new_n1888_), .A2(new_n1892_), .A3(new_n1894_), .ZN(new_n1895_));
  NOR2_X1   g1703(.A1(new_n1890_), .A2(new_n1891_), .ZN(new_n1896_));
  AOI221_X4 g1704(.A(new_n1887_), .B1(new_n1694_), .B2(new_n1698_), .C1(new_n1889_), .C2(new_n1699_), .ZN(new_n1897_));
  OAI21_X1  g1705(.A(new_n1893_), .B1(new_n1896_), .B2(new_n1897_), .ZN(new_n1898_));
  NAND3_X1  g1706(.A1(new_n1869_), .A2(new_n1895_), .A3(new_n1898_), .ZN(new_n1899_));
  NAND2_X1  g1707(.A1(new_n1898_), .A2(new_n1895_), .ZN(new_n1900_));
  NAND3_X1  g1708(.A1(new_n1900_), .A2(new_n1709_), .A3(new_n1718_), .ZN(new_n1901_));
  NAND2_X1  g1709(.A1(G188gat), .A2(G375gat), .ZN(new_n1902_));
  NAND3_X1  g1710(.A1(new_n1899_), .A2(new_n1901_), .A3(new_n1902_), .ZN(new_n1903_));
  INV_X1    g1711(.A(new_n1903_), .ZN(new_n1904_));
  AOI21_X1  g1712(.A(new_n1902_), .B1(new_n1899_), .B2(new_n1901_), .ZN(new_n1905_));
  OAI211_X1 g1713(.A(new_n1719_), .B(new_n1722_), .C1(new_n1904_), .C2(new_n1905_), .ZN(new_n1906_));
  INV_X1    g1714(.A(new_n1905_), .ZN(new_n1907_));
  AOI21_X1  g1715(.A(KEYINPUT79), .B1(new_n1907_), .B2(new_n1903_), .ZN(new_n1908_));
  NAND2_X1  g1716(.A1(new_n1722_), .A2(new_n1719_), .ZN(new_n1909_));
  AND2_X1   g1717(.A1(new_n1899_), .A2(new_n1901_), .ZN(new_n1910_));
  NAND2_X1  g1718(.A1(new_n1910_), .A2(KEYINPUT79), .ZN(new_n1911_));
  NAND2_X1  g1719(.A1(new_n1909_), .A2(new_n1911_), .ZN(new_n1912_));
  OAI211_X1 g1720(.A(new_n1867_), .B(new_n1906_), .C1(new_n1908_), .C2(new_n1912_), .ZN(new_n1913_));
  INV_X1    g1721(.A(new_n1913_), .ZN(new_n1914_));
  AOI22_X1  g1722(.A1(new_n1719_), .A2(new_n1722_), .B1(new_n1910_), .B2(KEYINPUT79), .ZN(new_n1915_));
  INV_X1    g1723(.A(KEYINPUT79), .ZN(new_n1916_));
  OAI21_X1  g1724(.A(new_n1916_), .B1(new_n1904_), .B2(new_n1905_), .ZN(new_n1917_));
  NAND2_X1  g1725(.A1(new_n1915_), .A2(new_n1917_), .ZN(new_n1918_));
  AOI21_X1  g1726(.A(new_n1867_), .B1(new_n1918_), .B2(new_n1906_), .ZN(new_n1919_));
  OAI21_X1  g1727(.A(new_n1865_), .B1(new_n1914_), .B2(new_n1919_), .ZN(new_n1920_));
  OAI21_X1  g1728(.A(new_n1906_), .B1(new_n1908_), .B2(new_n1912_), .ZN(new_n1921_));
  NAND2_X1  g1729(.A1(new_n1921_), .A2(new_n1866_), .ZN(new_n1922_));
  NAND2_X1  g1730(.A1(new_n1732_), .A2(new_n1729_), .ZN(new_n1923_));
  NAND3_X1  g1731(.A1(new_n1922_), .A2(new_n1923_), .A3(new_n1913_), .ZN(new_n1924_));
  NOR2_X1   g1732(.A1(new_n960_), .A2(new_n613_), .ZN(new_n1925_));
  NAND3_X1  g1733(.A1(new_n1920_), .A2(new_n1924_), .A3(new_n1925_), .ZN(new_n1926_));
  AOI21_X1  g1734(.A(new_n1925_), .B1(new_n1920_), .B2(new_n1924_), .ZN(new_n1927_));
  OAI21_X1  g1735(.A(new_n1926_), .B1(new_n1927_), .B2(KEYINPUT80), .ZN(new_n1928_));
  INV_X1    g1736(.A(KEYINPUT80), .ZN(new_n1929_));
  AOI211_X1 g1737(.A(new_n1929_), .B(new_n1925_), .C1(new_n1920_), .C2(new_n1924_), .ZN(new_n1930_));
  OAI21_X1  g1738(.A(new_n1864_), .B1(new_n1928_), .B2(new_n1930_), .ZN(new_n1931_));
  INV_X1    g1739(.A(new_n1927_), .ZN(new_n1932_));
  NAND3_X1  g1740(.A1(new_n1932_), .A2(new_n1863_), .A3(new_n1926_), .ZN(new_n1933_));
  AOI21_X1  g1741(.A(new_n1857_), .B1(new_n1931_), .B2(new_n1933_), .ZN(new_n1934_));
  INV_X1    g1742(.A(new_n1934_), .ZN(new_n1935_));
  NAND3_X1  g1743(.A1(new_n1931_), .A2(new_n1857_), .A3(new_n1933_), .ZN(new_n1936_));
  NAND2_X1  g1744(.A1(new_n1935_), .A2(new_n1936_), .ZN(new_n1937_));
  INV_X1    g1745(.A(new_n1937_), .ZN(new_n1938_));
  NAND2_X1  g1746(.A1(new_n1856_), .A2(new_n1938_), .ZN(new_n1939_));
  NAND2_X1  g1747(.A1(new_n1852_), .A2(new_n1850_), .ZN(new_n1940_));
  INV_X1    g1748(.A(new_n1940_), .ZN(new_n1941_));
  AOI21_X1  g1749(.A(KEYINPUT81), .B1(new_n1935_), .B2(new_n1936_), .ZN(new_n1942_));
  INV_X1    g1750(.A(KEYINPUT81), .ZN(new_n1943_));
  NOR2_X1   g1751(.A1(new_n1934_), .A2(new_n1943_), .ZN(new_n1944_));
  OAI21_X1  g1752(.A(new_n1941_), .B1(new_n1942_), .B2(new_n1944_), .ZN(new_n1945_));
  NOR2_X1   g1753(.A1(new_n532_), .A2(new_n768_), .ZN(new_n1946_));
  NAND3_X1  g1754(.A1(new_n1939_), .A2(new_n1945_), .A3(new_n1946_), .ZN(new_n1947_));
  INV_X1    g1755(.A(new_n1946_), .ZN(new_n1948_));
  AOI21_X1  g1756(.A(new_n1937_), .B1(new_n1853_), .B2(new_n1855_), .ZN(new_n1949_));
  INV_X1    g1757(.A(new_n1944_), .ZN(new_n1950_));
  AND3_X1   g1758(.A1(new_n1931_), .A2(new_n1857_), .A3(new_n1933_), .ZN(new_n1951_));
  OAI21_X1  g1759(.A(new_n1943_), .B1(new_n1951_), .B2(new_n1934_), .ZN(new_n1952_));
  AOI21_X1  g1760(.A(new_n1940_), .B1(new_n1950_), .B2(new_n1952_), .ZN(new_n1953_));
  OAI21_X1  g1761(.A(new_n1948_), .B1(new_n1949_), .B2(new_n1953_), .ZN(new_n1954_));
  NAND2_X1  g1762(.A1(new_n1774_), .A2(KEYINPUT77), .ZN(new_n1955_));
  INV_X1    g1763(.A(KEYINPUT77), .ZN(new_n1956_));
  NAND3_X1  g1764(.A1(new_n1757_), .A2(new_n1956_), .A3(new_n1761_), .ZN(new_n1957_));
  NAND3_X1  g1765(.A1(new_n1955_), .A2(new_n1771_), .A3(new_n1957_), .ZN(new_n1958_));
  NAND2_X1  g1766(.A1(new_n1958_), .A2(KEYINPUT76), .ZN(new_n1959_));
  NAND3_X1  g1767(.A1(new_n1947_), .A2(new_n1954_), .A3(new_n1959_), .ZN(new_n1960_));
  AND2_X1   g1768(.A1(new_n1789_), .A2(new_n1958_), .ZN(new_n1961_));
  NAND2_X1  g1769(.A1(new_n1960_), .A2(new_n1961_), .ZN(new_n1962_));
  NOR2_X1   g1770(.A1(new_n452_), .A2(new_n918_), .ZN(new_n1963_));
  INV_X1    g1771(.A(new_n1963_), .ZN(new_n1964_));
  NAND2_X1  g1772(.A1(new_n1789_), .A2(new_n1958_), .ZN(new_n1965_));
  NAND4_X1  g1773(.A1(new_n1965_), .A2(new_n1954_), .A3(new_n1947_), .A4(new_n1959_), .ZN(new_n1966_));
  AND3_X1   g1774(.A1(new_n1962_), .A2(new_n1964_), .A3(new_n1966_), .ZN(new_n1967_));
  AOI21_X1  g1775(.A(new_n1964_), .B1(new_n1962_), .B2(new_n1966_), .ZN(new_n1968_));
  OAI21_X1  g1776(.A(new_n1848_), .B1(new_n1967_), .B2(new_n1968_), .ZN(new_n1969_));
  NAND2_X1  g1777(.A1(new_n1962_), .A2(new_n1966_), .ZN(new_n1970_));
  NAND2_X1  g1778(.A1(new_n1970_), .A2(new_n1963_), .ZN(new_n1971_));
  NAND2_X1  g1779(.A1(new_n1791_), .A2(new_n1790_), .ZN(new_n1972_));
  NAND3_X1  g1780(.A1(new_n1962_), .A2(new_n1964_), .A3(new_n1966_), .ZN(new_n1973_));
  NAND3_X1  g1781(.A1(new_n1971_), .A2(new_n1972_), .A3(new_n1973_), .ZN(new_n1974_));
  NOR2_X1   g1782(.A1(new_n310_), .A2(new_n1419_), .ZN(new_n1975_));
  INV_X1    g1783(.A(new_n1975_), .ZN(new_n1976_));
  AND3_X1   g1784(.A1(new_n1969_), .A2(new_n1974_), .A3(new_n1976_), .ZN(new_n1977_));
  AOI21_X1  g1785(.A(new_n1976_), .B1(new_n1969_), .B2(new_n1974_), .ZN(new_n1978_));
  OAI211_X1 g1786(.A(new_n1794_), .B(new_n1805_), .C1(new_n1977_), .C2(new_n1978_), .ZN(new_n1979_));
  NOR2_X1   g1787(.A1(new_n241_), .A2(new_n1426_), .ZN(new_n1980_));
  INV_X1    g1788(.A(new_n1980_), .ZN(new_n1981_));
  NOR3_X1   g1789(.A1(new_n1967_), .A2(new_n1968_), .A3(new_n1848_), .ZN(new_n1982_));
  AOI21_X1  g1790(.A(new_n1972_), .B1(new_n1971_), .B2(new_n1973_), .ZN(new_n1983_));
  OAI21_X1  g1791(.A(new_n1975_), .B1(new_n1982_), .B2(new_n1983_), .ZN(new_n1984_));
  AOI21_X1  g1792(.A(new_n1663_), .B1(new_n1791_), .B2(new_n1793_), .ZN(new_n1985_));
  OAI21_X1  g1793(.A(new_n1794_), .B1(new_n1985_), .B2(new_n1795_), .ZN(new_n1986_));
  NAND3_X1  g1794(.A1(new_n1969_), .A2(new_n1974_), .A3(new_n1976_), .ZN(new_n1987_));
  NAND3_X1  g1795(.A1(new_n1984_), .A2(new_n1986_), .A3(new_n1987_), .ZN(new_n1988_));
  NAND3_X1  g1796(.A1(new_n1979_), .A2(new_n1981_), .A3(new_n1988_), .ZN(new_n1989_));
  AND3_X1   g1797(.A1(new_n1984_), .A2(new_n1986_), .A3(new_n1987_), .ZN(new_n1990_));
  AOI21_X1  g1798(.A(new_n1986_), .B1(new_n1984_), .B2(new_n1987_), .ZN(new_n1991_));
  OAI21_X1  g1799(.A(new_n1980_), .B1(new_n1990_), .B2(new_n1991_), .ZN(new_n1992_));
  NAND3_X1  g1800(.A1(new_n1846_), .A2(new_n1989_), .A3(new_n1992_), .ZN(new_n1993_));
  NAND2_X1  g1801(.A1(new_n1845_), .A2(new_n1806_), .ZN(new_n1994_));
  INV_X1    g1802(.A(new_n1994_), .ZN(new_n1995_));
  NAND2_X1  g1803(.A1(new_n1993_), .A2(new_n1995_), .ZN(new_n1996_));
  NOR2_X1   g1804(.A1(new_n215_), .A2(new_n1438_), .ZN(new_n1997_));
  INV_X1    g1805(.A(new_n1997_), .ZN(new_n1998_));
  NAND4_X1  g1806(.A1(new_n1994_), .A2(new_n1846_), .A3(new_n1989_), .A4(new_n1992_), .ZN(new_n1999_));
  AND3_X1   g1807(.A1(new_n1996_), .A2(new_n1998_), .A3(new_n1999_), .ZN(new_n2000_));
  AOI21_X1  g1808(.A(new_n1998_), .B1(new_n1996_), .B2(new_n1999_), .ZN(new_n2001_));
  OAI211_X1 g1809(.A(new_n1828_), .B(new_n1844_), .C1(new_n2000_), .C2(new_n2001_), .ZN(new_n2002_));
  NAND2_X1  g1810(.A1(new_n1828_), .A2(new_n1844_), .ZN(new_n2003_));
  NAND3_X1  g1811(.A1(new_n1996_), .A2(new_n1998_), .A3(new_n1999_), .ZN(new_n2004_));
  NOR3_X1   g1812(.A1(new_n1990_), .A2(new_n1991_), .A3(new_n1980_), .ZN(new_n2005_));
  AOI21_X1  g1813(.A(new_n1981_), .B1(new_n1979_), .B2(new_n1988_), .ZN(new_n2006_));
  NOR2_X1   g1814(.A1(new_n2005_), .A2(new_n2006_), .ZN(new_n2007_));
  AOI21_X1  g1815(.A(new_n1994_), .B1(new_n2007_), .B2(new_n1846_), .ZN(new_n2008_));
  INV_X1    g1816(.A(new_n1999_), .ZN(new_n2009_));
  OAI21_X1  g1817(.A(new_n1997_), .B1(new_n2008_), .B2(new_n2009_), .ZN(new_n2010_));
  NAND3_X1  g1818(.A1(new_n2003_), .A2(new_n2004_), .A3(new_n2010_), .ZN(new_n2011_));
  NOR2_X1   g1819(.A1(new_n205_), .A2(new_n1654_), .ZN(new_n2012_));
  XOR2_X1   g1820(.A(new_n2012_), .B(KEYINPUT83), .Z(new_n2013_));
  AND3_X1   g1821(.A1(new_n2002_), .A2(new_n2011_), .A3(new_n2013_), .ZN(new_n2014_));
  AOI21_X1  g1822(.A(new_n2013_), .B1(new_n2002_), .B2(new_n2011_), .ZN(new_n2015_));
  OAI21_X1  g1823(.A(new_n1843_), .B1(new_n2014_), .B2(new_n2015_), .ZN(new_n2016_));
  NAND2_X1  g1824(.A1(new_n2002_), .A2(new_n2011_), .ZN(new_n2017_));
  INV_X1    g1825(.A(new_n2013_), .ZN(new_n2018_));
  NAND2_X1  g1826(.A1(new_n2017_), .A2(new_n2018_), .ZN(new_n2019_));
  OAI21_X1  g1827(.A(new_n1837_), .B1(new_n1830_), .B2(new_n1831_), .ZN(new_n2020_));
  NAND3_X1  g1828(.A1(new_n2002_), .A2(new_n2011_), .A3(new_n2012_), .ZN(new_n2021_));
  NAND3_X1  g1829(.A1(new_n2019_), .A2(new_n2020_), .A3(new_n2021_), .ZN(new_n2022_));
  NAND2_X1  g1830(.A1(new_n2016_), .A2(new_n2022_), .ZN(new_n2023_));
  XNOR2_X1  g1831(.A(new_n2023_), .B(new_n1839_), .ZN(G6160gat));
  OAI21_X1  g1832(.A(new_n1988_), .B1(new_n1991_), .B2(new_n1980_), .ZN(new_n2025_));
  INV_X1    g1833(.A(new_n2025_), .ZN(new_n2026_));
  AOI21_X1  g1834(.A(new_n1982_), .B1(new_n1976_), .B2(new_n1969_), .ZN(new_n2027_));
  NAND3_X1  g1835(.A1(new_n1965_), .A2(new_n1954_), .A3(new_n1947_), .ZN(new_n2028_));
  AND2_X1   g1836(.A1(new_n1973_), .A2(new_n2028_), .ZN(new_n2029_));
  INV_X1    g1837(.A(KEYINPUT87), .ZN(new_n2030_));
  NAND2_X1  g1838(.A1(new_n2028_), .A2(new_n2030_), .ZN(new_n2031_));
  NAND2_X1  g1839(.A1(new_n1931_), .A2(new_n1857_), .ZN(new_n2032_));
  NAND2_X1  g1840(.A1(new_n2032_), .A2(new_n1933_), .ZN(new_n2033_));
  INV_X1    g1841(.A(KEYINPUT86), .ZN(new_n2034_));
  OR2_X1    g1842(.A1(new_n1924_), .A2(new_n2034_), .ZN(new_n2035_));
  INV_X1    g1843(.A(new_n1925_), .ZN(new_n2036_));
  NAND3_X1  g1844(.A1(new_n1920_), .A2(new_n1924_), .A3(new_n2036_), .ZN(new_n2037_));
  NAND2_X1  g1845(.A1(new_n1924_), .A2(new_n2034_), .ZN(new_n2038_));
  NAND3_X1  g1846(.A1(new_n2035_), .A2(new_n2037_), .A3(new_n2038_), .ZN(new_n2039_));
  OAI21_X1  g1847(.A(new_n1888_), .B1(new_n1897_), .B2(new_n1893_), .ZN(new_n2040_));
  INV_X1    g1848(.A(new_n1886_), .ZN(new_n2041_));
  NOR2_X1   g1849(.A1(new_n2041_), .A2(new_n1885_), .ZN(new_n2042_));
  NAND3_X1  g1850(.A1(new_n1874_), .A2(new_n1877_), .A3(new_n1875_), .ZN(new_n2043_));
  NAND2_X1  g1851(.A1(new_n2043_), .A2(new_n1874_), .ZN(new_n2044_));
  OAI21_X1  g1852(.A(new_n2044_), .B1(new_n1872_), .B2(new_n232_), .ZN(new_n2045_));
  NAND3_X1  g1853(.A1(new_n2043_), .A2(G324gat), .A3(new_n1874_), .ZN(new_n2046_));
  NAND2_X1  g1854(.A1(new_n2045_), .A2(new_n2046_), .ZN(new_n2047_));
  NAND2_X1  g1855(.A1(G239gat), .A2(G341gat), .ZN(new_n2048_));
  XOR2_X1   g1856(.A(new_n2047_), .B(new_n2048_), .Z(new_n2049_));
  NAND2_X1  g1857(.A1(new_n2042_), .A2(new_n2049_), .ZN(new_n2050_));
  NOR2_X1   g1858(.A1(new_n1882_), .A2(new_n1883_), .ZN(new_n2051_));
  NOR2_X1   g1859(.A1(new_n2051_), .A2(new_n2041_), .ZN(new_n2052_));
  OAI21_X1  g1860(.A(new_n2050_), .B1(new_n2052_), .B2(new_n2049_), .ZN(new_n2053_));
  NOR2_X1   g1861(.A1(new_n300_), .A2(new_n1681_), .ZN(new_n2054_));
  NAND2_X1  g1862(.A1(new_n2053_), .A2(new_n2054_), .ZN(new_n2055_));
  OAI221_X1 g1863(.A(new_n2050_), .B1(new_n1681_), .B2(new_n300_), .C1(new_n2052_), .C2(new_n2049_), .ZN(new_n2056_));
  NAND3_X1  g1864(.A1(new_n2040_), .A2(new_n2055_), .A3(new_n2056_), .ZN(new_n2057_));
  NAND2_X1  g1865(.A1(new_n2055_), .A2(new_n2056_), .ZN(new_n2058_));
  NAND3_X1  g1866(.A1(new_n1895_), .A2(new_n1888_), .A3(new_n2058_), .ZN(new_n2059_));
  NAND2_X1  g1867(.A1(new_n2057_), .A2(new_n2059_), .ZN(new_n2060_));
  NOR2_X1   g1868(.A1(new_n944_), .A2(new_n355_), .ZN(new_n2061_));
  NAND2_X1  g1869(.A1(new_n2060_), .A2(new_n2061_), .ZN(new_n2062_));
  INV_X1    g1870(.A(new_n2061_), .ZN(new_n2063_));
  NAND3_X1  g1871(.A1(new_n2057_), .A2(new_n2059_), .A3(new_n2063_), .ZN(new_n2064_));
  NAND2_X1  g1872(.A1(new_n2062_), .A2(new_n2064_), .ZN(new_n2065_));
  NAND2_X1  g1873(.A1(new_n2065_), .A2(KEYINPUT84), .ZN(new_n2066_));
  NAND2_X1  g1874(.A1(new_n1903_), .A2(new_n1899_), .ZN(new_n2067_));
  INV_X1    g1875(.A(KEYINPUT84), .ZN(new_n2068_));
  NAND3_X1  g1876(.A1(new_n2062_), .A2(new_n2068_), .A3(new_n2064_), .ZN(new_n2069_));
  NAND3_X1  g1877(.A1(new_n2066_), .A2(new_n2067_), .A3(new_n2069_), .ZN(new_n2070_));
  NAND4_X1  g1878(.A1(new_n2065_), .A2(KEYINPUT84), .A3(new_n1903_), .A4(new_n1899_), .ZN(new_n2071_));
  NAND2_X1  g1879(.A1(new_n2070_), .A2(new_n2071_), .ZN(new_n2072_));
  NOR2_X1   g1880(.A1(new_n1093_), .A2(new_n601_), .ZN(new_n2073_));
  INV_X1    g1881(.A(new_n2073_), .ZN(new_n2074_));
  NOR2_X1   g1882(.A1(new_n2074_), .A2(KEYINPUT85), .ZN(new_n2075_));
  INV_X1    g1883(.A(new_n2075_), .ZN(new_n2076_));
  NAND2_X1  g1884(.A1(new_n2072_), .A2(new_n2076_), .ZN(new_n2077_));
  XOR2_X1   g1885(.A(new_n2073_), .B(KEYINPUT85), .Z(new_n2078_));
  NAND3_X1  g1886(.A1(new_n2070_), .A2(new_n2071_), .A3(new_n2078_), .ZN(new_n2079_));
  NAND4_X1  g1887(.A1(new_n2077_), .A2(new_n1913_), .A3(new_n1918_), .A4(new_n2079_), .ZN(new_n2080_));
  AOI21_X1  g1888(.A(new_n1909_), .B1(new_n1903_), .B2(new_n1907_), .ZN(new_n2081_));
  OAI21_X1  g1889(.A(new_n1918_), .B1(new_n2081_), .B2(new_n1866_), .ZN(new_n2082_));
  AND3_X1   g1890(.A1(new_n2070_), .A2(new_n2071_), .A3(new_n2078_), .ZN(new_n2083_));
  AOI21_X1  g1891(.A(new_n2075_), .B1(new_n2070_), .B2(new_n2071_), .ZN(new_n2084_));
  OAI21_X1  g1892(.A(new_n2082_), .B1(new_n2083_), .B2(new_n2084_), .ZN(new_n2085_));
  NAND2_X1  g1893(.A1(G171gat), .A2(G409gat), .ZN(new_n2086_));
  AND3_X1   g1894(.A1(new_n2080_), .A2(new_n2085_), .A3(new_n2086_), .ZN(new_n2087_));
  AOI21_X1  g1895(.A(new_n2086_), .B1(new_n2080_), .B2(new_n2085_), .ZN(new_n2088_));
  NOR2_X1   g1896(.A1(new_n2087_), .A2(new_n2088_), .ZN(new_n2089_));
  OR2_X1    g1897(.A1(new_n2039_), .A2(new_n2089_), .ZN(new_n2090_));
  NAND2_X1  g1898(.A1(G154gat), .A2(G426gat), .ZN(new_n2091_));
  NAND2_X1  g1899(.A1(new_n2039_), .A2(new_n2089_), .ZN(new_n2092_));
  AND3_X1   g1900(.A1(new_n2090_), .A2(new_n2091_), .A3(new_n2092_), .ZN(new_n2093_));
  AOI21_X1  g1901(.A(new_n2091_), .B1(new_n2090_), .B2(new_n2092_), .ZN(new_n2094_));
  OAI21_X1  g1902(.A(new_n2033_), .B1(new_n2093_), .B2(new_n2094_), .ZN(new_n2095_));
  AND2_X1   g1903(.A1(new_n2039_), .A2(new_n2089_), .ZN(new_n2096_));
  NOR2_X1   g1904(.A1(new_n2039_), .A2(new_n2089_), .ZN(new_n2097_));
  OAI211_X1 g1905(.A(G154gat), .B(G426gat), .C1(new_n2096_), .C2(new_n2097_), .ZN(new_n2098_));
  NAND3_X1  g1906(.A1(new_n2090_), .A2(new_n2091_), .A3(new_n2092_), .ZN(new_n2099_));
  NAND4_X1  g1907(.A1(new_n2098_), .A2(new_n2099_), .A3(new_n1933_), .A4(new_n2032_), .ZN(new_n2100_));
  NAND2_X1  g1908(.A1(new_n2095_), .A2(new_n2100_), .ZN(new_n2101_));
  NAND3_X1  g1909(.A1(new_n2101_), .A2(G137gat), .A3(G443gat), .ZN(new_n2102_));
  OAI211_X1 g1910(.A(new_n2095_), .B(new_n2100_), .C1(new_n651_), .C2(new_n768_), .ZN(new_n2103_));
  NAND2_X1  g1911(.A1(new_n2102_), .A2(new_n2103_), .ZN(new_n2104_));
  NAND2_X1  g1912(.A1(new_n1950_), .A2(new_n1952_), .ZN(new_n2105_));
  NAND2_X1  g1913(.A1(new_n1856_), .A2(new_n2105_), .ZN(new_n2106_));
  AND3_X1   g1914(.A1(new_n1954_), .A2(new_n2104_), .A3(new_n2106_), .ZN(new_n2107_));
  AOI21_X1  g1915(.A(new_n2104_), .B1(new_n1954_), .B2(new_n2106_), .ZN(new_n2108_));
  NOR2_X1   g1916(.A1(new_n532_), .A2(new_n918_), .ZN(new_n2109_));
  NOR3_X1   g1917(.A1(new_n2107_), .A2(new_n2108_), .A3(new_n2109_), .ZN(new_n2110_));
  INV_X1    g1918(.A(new_n2109_), .ZN(new_n2111_));
  AND2_X1   g1919(.A1(new_n2102_), .A2(new_n2103_), .ZN(new_n2112_));
  AOI21_X1  g1920(.A(new_n1946_), .B1(new_n1939_), .B2(new_n1945_), .ZN(new_n2113_));
  INV_X1    g1921(.A(new_n2106_), .ZN(new_n2114_));
  OAI21_X1  g1922(.A(new_n2112_), .B1(new_n2113_), .B2(new_n2114_), .ZN(new_n2115_));
  NAND3_X1  g1923(.A1(new_n1954_), .A2(new_n2104_), .A3(new_n2106_), .ZN(new_n2116_));
  AOI21_X1  g1924(.A(new_n2111_), .B1(new_n2115_), .B2(new_n2116_), .ZN(new_n2117_));
  OAI21_X1  g1925(.A(new_n2031_), .B1(new_n2110_), .B2(new_n2117_), .ZN(new_n2118_));
  NAND2_X1  g1926(.A1(new_n2029_), .A2(new_n2118_), .ZN(new_n2119_));
  NOR2_X1   g1927(.A1(new_n452_), .A2(new_n1419_), .ZN(new_n2120_));
  OAI21_X1  g1928(.A(new_n2109_), .B1(new_n2107_), .B2(new_n2108_), .ZN(new_n2121_));
  NAND3_X1  g1929(.A1(new_n2115_), .A2(new_n2111_), .A3(new_n2116_), .ZN(new_n2122_));
  AOI22_X1  g1930(.A1(new_n2121_), .A2(new_n2122_), .B1(new_n2030_), .B2(new_n2028_), .ZN(new_n2123_));
  NAND2_X1  g1931(.A1(new_n1973_), .A2(new_n2028_), .ZN(new_n2124_));
  NAND2_X1  g1932(.A1(new_n2123_), .A2(new_n2124_), .ZN(new_n2125_));
  AND3_X1   g1933(.A1(new_n2119_), .A2(new_n2120_), .A3(new_n2125_), .ZN(new_n2126_));
  AOI21_X1  g1934(.A(new_n2120_), .B1(new_n2119_), .B2(new_n2125_), .ZN(new_n2127_));
  OAI21_X1  g1935(.A(new_n2027_), .B1(new_n2126_), .B2(new_n2127_), .ZN(new_n2128_));
  NOR2_X1   g1936(.A1(new_n2029_), .A2(new_n2118_), .ZN(new_n2129_));
  NOR2_X1   g1937(.A1(new_n2123_), .A2(new_n2124_), .ZN(new_n2130_));
  OAI22_X1  g1938(.A1(new_n2129_), .A2(new_n2130_), .B1(new_n452_), .B2(new_n1419_), .ZN(new_n2131_));
  NAND2_X1  g1939(.A1(new_n1987_), .A2(new_n1974_), .ZN(new_n2132_));
  NAND3_X1  g1940(.A1(new_n2119_), .A2(new_n2120_), .A3(new_n2125_), .ZN(new_n2133_));
  NAND3_X1  g1941(.A1(new_n2131_), .A2(new_n2132_), .A3(new_n2133_), .ZN(new_n2134_));
  NOR2_X1   g1942(.A1(new_n310_), .A2(new_n1426_), .ZN(new_n2135_));
  INV_X1    g1943(.A(new_n2135_), .ZN(new_n2136_));
  AND3_X1   g1944(.A1(new_n2128_), .A2(new_n2134_), .A3(new_n2136_), .ZN(new_n2137_));
  AOI21_X1  g1945(.A(new_n2136_), .B1(new_n2128_), .B2(new_n2134_), .ZN(new_n2138_));
  OAI21_X1  g1946(.A(new_n2026_), .B1(new_n2137_), .B2(new_n2138_), .ZN(new_n2139_));
  NOR3_X1   g1947(.A1(new_n2126_), .A2(new_n2127_), .A3(new_n2027_), .ZN(new_n2140_));
  AOI21_X1  g1948(.A(new_n2132_), .B1(new_n2131_), .B2(new_n2133_), .ZN(new_n2141_));
  OAI21_X1  g1949(.A(new_n2135_), .B1(new_n2140_), .B2(new_n2141_), .ZN(new_n2142_));
  NAND3_X1  g1950(.A1(new_n2128_), .A2(new_n2134_), .A3(new_n2136_), .ZN(new_n2143_));
  NAND3_X1  g1951(.A1(new_n2142_), .A2(new_n2025_), .A3(new_n2143_), .ZN(new_n2144_));
  NAND2_X1  g1952(.A1(G69gat), .A2(G511gat), .ZN(new_n2145_));
  AND3_X1   g1953(.A1(new_n2139_), .A2(new_n2144_), .A3(new_n2145_), .ZN(new_n2146_));
  AOI21_X1  g1954(.A(new_n2145_), .B1(new_n2139_), .B2(new_n2144_), .ZN(new_n2147_));
  NOR2_X1   g1955(.A1(new_n2146_), .A2(new_n2147_), .ZN(new_n2148_));
  NAND2_X1  g1956(.A1(new_n2007_), .A2(new_n1994_), .ZN(new_n2149_));
  NAND2_X1  g1957(.A1(new_n2004_), .A2(new_n2149_), .ZN(new_n2150_));
  NAND2_X1  g1958(.A1(new_n2148_), .A2(new_n2150_), .ZN(new_n2151_));
  OAI211_X1 g1959(.A(new_n2004_), .B(new_n2149_), .C1(new_n2146_), .C2(new_n2147_), .ZN(new_n2152_));
  NAND2_X1  g1960(.A1(new_n2151_), .A2(new_n2152_), .ZN(new_n2153_));
  NOR2_X1   g1961(.A1(new_n215_), .A2(new_n1654_), .ZN(new_n2154_));
  NAND2_X1  g1962(.A1(new_n2153_), .A2(new_n2154_), .ZN(new_n2155_));
  INV_X1    g1963(.A(new_n2154_), .ZN(new_n2156_));
  NAND3_X1  g1964(.A1(new_n2151_), .A2(new_n2156_), .A3(new_n2152_), .ZN(new_n2157_));
  NAND2_X1  g1965(.A1(new_n2155_), .A2(new_n2157_), .ZN(new_n2158_));
  INV_X1    g1966(.A(new_n2012_), .ZN(new_n2159_));
  NAND2_X1  g1967(.A1(new_n2002_), .A2(new_n2159_), .ZN(new_n2160_));
  NAND2_X1  g1968(.A1(new_n2160_), .A2(new_n2011_), .ZN(new_n2161_));
  INV_X1    g1969(.A(new_n2161_), .ZN(new_n2162_));
  AOI21_X1  g1970(.A(KEYINPUT88), .B1(new_n2158_), .B2(new_n2162_), .ZN(new_n2163_));
  NAND2_X1  g1971(.A1(new_n2011_), .A2(new_n2013_), .ZN(new_n2164_));
  NAND4_X1  g1972(.A1(new_n2155_), .A2(new_n2002_), .A3(new_n2157_), .A4(new_n2164_), .ZN(new_n2165_));
  INV_X1    g1973(.A(new_n2157_), .ZN(new_n2166_));
  AOI21_X1  g1974(.A(new_n2156_), .B1(new_n2151_), .B2(new_n2152_), .ZN(new_n2167_));
  OAI21_X1  g1975(.A(new_n2161_), .B1(new_n2166_), .B2(new_n2167_), .ZN(new_n2168_));
  AOI22_X1  g1976(.A1(new_n2163_), .A2(new_n2165_), .B1(KEYINPUT88), .B2(new_n2168_), .ZN(new_n2169_));
  NAND3_X1  g1977(.A1(new_n2002_), .A2(new_n2011_), .A3(new_n2013_), .ZN(new_n2170_));
  AOI21_X1  g1978(.A(new_n1843_), .B1(new_n2019_), .B2(new_n2170_), .ZN(new_n2171_));
  AOI21_X1  g1979(.A(new_n2171_), .B1(new_n2023_), .B2(new_n1839_), .ZN(new_n2172_));
  XNOR2_X1  g1980(.A(new_n2169_), .B(new_n2172_), .ZN(G6170gat));
  OAI21_X1  g1981(.A(new_n2165_), .B1(new_n2169_), .B2(new_n2172_), .ZN(new_n2174_));
  NOR2_X1   g1982(.A1(new_n241_), .A2(new_n1654_), .ZN(new_n2175_));
  NOR2_X1   g1983(.A1(new_n2137_), .A2(new_n2140_), .ZN(new_n2176_));
  INV_X1    g1984(.A(new_n2176_), .ZN(new_n2177_));
  NOR2_X1   g1985(.A1(new_n651_), .A2(new_n918_), .ZN(new_n2178_));
  NOR2_X1   g1986(.A1(new_n960_), .A2(new_n768_), .ZN(new_n2179_));
  INV_X1    g1987(.A(new_n2179_), .ZN(new_n2180_));
  XNOR2_X1  g1988(.A(new_n2096_), .B(KEYINPUT89), .ZN(new_n2181_));
  NOR2_X1   g1989(.A1(new_n2181_), .A2(new_n2093_), .ZN(new_n2182_));
  NAND3_X1  g1990(.A1(new_n2070_), .A2(new_n2071_), .A3(new_n2074_), .ZN(new_n2183_));
  NAND3_X1  g1991(.A1(new_n2067_), .A2(new_n2064_), .A3(new_n2062_), .ZN(new_n2184_));
  NAND2_X1  g1992(.A1(new_n2183_), .A2(new_n2184_), .ZN(new_n2185_));
  AND2_X1   g1993(.A1(new_n2064_), .A2(new_n2057_), .ZN(new_n2186_));
  NAND3_X1  g1994(.A1(new_n2045_), .A2(new_n2048_), .A3(new_n2046_), .ZN(new_n2187_));
  NAND2_X1  g1995(.A1(new_n2187_), .A2(new_n2045_), .ZN(new_n2188_));
  NAND2_X1  g1996(.A1(G256gat), .A2(G341gat), .ZN(new_n2189_));
  OR2_X1    g1997(.A1(new_n2188_), .A2(new_n2189_), .ZN(new_n2190_));
  NAND2_X1  g1998(.A1(new_n2188_), .A2(new_n2189_), .ZN(new_n2191_));
  NAND2_X1  g1999(.A1(new_n2190_), .A2(new_n2191_), .ZN(new_n2192_));
  NAND2_X1  g2000(.A1(new_n299_), .A2(G239gat), .ZN(new_n2193_));
  XNOR2_X1  g2001(.A(new_n2192_), .B(new_n2193_), .ZN(new_n2194_));
  OAI21_X1  g2002(.A(new_n2054_), .B1(new_n2042_), .B2(new_n2049_), .ZN(new_n2195_));
  NAND3_X1  g2003(.A1(new_n2194_), .A2(new_n2050_), .A3(new_n2195_), .ZN(new_n2196_));
  INV_X1    g2004(.A(new_n2196_), .ZN(new_n2197_));
  AOI21_X1  g2005(.A(new_n2194_), .B1(new_n2050_), .B2(new_n2195_), .ZN(new_n2198_));
  NOR2_X1   g2006(.A1(new_n2197_), .A2(new_n2198_), .ZN(new_n2199_));
  NAND2_X1  g2007(.A1(G222gat), .A2(G375gat), .ZN(new_n2200_));
  XNOR2_X1  g2008(.A(new_n2199_), .B(new_n2200_), .ZN(new_n2201_));
  OR2_X1    g2009(.A1(new_n2186_), .A2(new_n2201_), .ZN(new_n2202_));
  NAND2_X1  g2010(.A1(new_n2186_), .A2(new_n2201_), .ZN(new_n2203_));
  OAI211_X1 g2011(.A(new_n2202_), .B(new_n2203_), .C1(new_n944_), .C2(new_n601_), .ZN(new_n2204_));
  NAND2_X1  g2012(.A1(new_n2202_), .A2(new_n2203_), .ZN(new_n2205_));
  NAND3_X1  g2013(.A1(new_n2205_), .A2(G205gat), .A3(G392gat), .ZN(new_n2206_));
  AND3_X1   g2014(.A1(new_n2185_), .A2(new_n2204_), .A3(new_n2206_), .ZN(new_n2207_));
  AOI21_X1  g2015(.A(new_n2185_), .B1(new_n2204_), .B2(new_n2206_), .ZN(new_n2208_));
  NOR2_X1   g2016(.A1(new_n1093_), .A2(new_n613_), .ZN(new_n2209_));
  OR3_X1    g2017(.A1(new_n2207_), .A2(new_n2208_), .A3(new_n2209_), .ZN(new_n2210_));
  NAND3_X1  g2018(.A1(new_n2080_), .A2(new_n2085_), .A3(new_n2086_), .ZN(new_n2211_));
  NAND2_X1  g2019(.A1(new_n2211_), .A2(new_n2085_), .ZN(new_n2212_));
  OAI21_X1  g2020(.A(new_n2209_), .B1(new_n2207_), .B2(new_n2208_), .ZN(new_n2213_));
  NAND3_X1  g2021(.A1(new_n2210_), .A2(new_n2212_), .A3(new_n2213_), .ZN(new_n2214_));
  INV_X1    g2022(.A(new_n2214_), .ZN(new_n2215_));
  NOR2_X1   g2023(.A1(new_n799_), .A2(new_n624_), .ZN(new_n2216_));
  AOI21_X1  g2024(.A(new_n2212_), .B1(new_n2210_), .B2(new_n2213_), .ZN(new_n2217_));
  NOR3_X1   g2025(.A1(new_n2215_), .A2(new_n2216_), .A3(new_n2217_), .ZN(new_n2218_));
  INV_X1    g2026(.A(new_n2218_), .ZN(new_n2219_));
  OAI21_X1  g2027(.A(new_n2216_), .B1(new_n2215_), .B2(new_n2217_), .ZN(new_n2220_));
  NAND2_X1  g2028(.A1(new_n2219_), .A2(new_n2220_), .ZN(new_n2221_));
  OR2_X1    g2029(.A1(new_n2182_), .A2(new_n2221_), .ZN(new_n2222_));
  NAND2_X1  g2030(.A1(new_n2182_), .A2(new_n2221_), .ZN(new_n2223_));
  AOI21_X1  g2031(.A(new_n2180_), .B1(new_n2222_), .B2(new_n2223_), .ZN(new_n2224_));
  INV_X1    g2032(.A(new_n2224_), .ZN(new_n2225_));
  NAND2_X1  g2033(.A1(new_n2103_), .A2(new_n2100_), .ZN(new_n2226_));
  NAND3_X1  g2034(.A1(new_n2222_), .A2(new_n2180_), .A3(new_n2223_), .ZN(new_n2227_));
  AND3_X1   g2035(.A1(new_n2225_), .A2(new_n2226_), .A3(new_n2227_), .ZN(new_n2228_));
  AOI21_X1  g2036(.A(new_n2226_), .B1(new_n2225_), .B2(new_n2227_), .ZN(new_n2229_));
  OAI21_X1  g2037(.A(new_n2178_), .B1(new_n2228_), .B2(new_n2229_), .ZN(new_n2230_));
  INV_X1    g2038(.A(new_n2227_), .ZN(new_n2231_));
  OAI211_X1 g2039(.A(new_n2100_), .B(new_n2103_), .C1(new_n2231_), .C2(new_n2224_), .ZN(new_n2232_));
  NAND3_X1  g2040(.A1(new_n2225_), .A2(new_n2226_), .A3(new_n2227_), .ZN(new_n2233_));
  OAI211_X1 g2041(.A(new_n2232_), .B(new_n2233_), .C1(new_n651_), .C2(new_n918_), .ZN(new_n2234_));
  NAND2_X1  g2042(.A1(new_n2230_), .A2(new_n2234_), .ZN(new_n2235_));
  NOR2_X1   g2043(.A1(new_n2110_), .A2(new_n2108_), .ZN(new_n2236_));
  OR2_X1    g2044(.A1(new_n2235_), .A2(new_n2236_), .ZN(new_n2237_));
  NAND2_X1  g2045(.A1(new_n2235_), .A2(new_n2236_), .ZN(new_n2238_));
  OAI21_X1  g2046(.A(KEYINPUT90), .B1(new_n532_), .B2(new_n1419_), .ZN(new_n2239_));
  AND3_X1   g2047(.A1(new_n2237_), .A2(new_n2238_), .A3(new_n2239_), .ZN(new_n2240_));
  OR3_X1    g2048(.A1(new_n532_), .A2(new_n1419_), .A3(KEYINPUT90), .ZN(new_n2241_));
  AOI22_X1  g2049(.A1(new_n2237_), .A2(new_n2238_), .B1(new_n2239_), .B2(new_n2241_), .ZN(new_n2242_));
  NOR2_X1   g2050(.A1(new_n2240_), .A2(new_n2242_), .ZN(new_n2243_));
  NOR3_X1   g2051(.A1(new_n2029_), .A2(new_n2110_), .A3(new_n2117_), .ZN(new_n2244_));
  NOR2_X1   g2052(.A1(new_n2127_), .A2(new_n2244_), .ZN(new_n2245_));
  OR2_X1    g2053(.A1(new_n2243_), .A2(new_n2245_), .ZN(new_n2246_));
  NAND2_X1  g2054(.A1(new_n2243_), .A2(new_n2245_), .ZN(new_n2247_));
  NAND2_X1  g2055(.A1(G103gat), .A2(G494gat), .ZN(new_n2248_));
  NAND2_X1  g2056(.A1(new_n2248_), .A2(KEYINPUT91), .ZN(new_n2249_));
  NAND3_X1  g2057(.A1(new_n2246_), .A2(new_n2247_), .A3(new_n2249_), .ZN(new_n2250_));
  INV_X1    g2058(.A(new_n2250_), .ZN(new_n2251_));
  OR2_X1    g2059(.A1(new_n2248_), .A2(KEYINPUT91), .ZN(new_n2252_));
  AOI22_X1  g2060(.A1(new_n2246_), .A2(new_n2247_), .B1(new_n2249_), .B2(new_n2252_), .ZN(new_n2253_));
  OAI21_X1  g2061(.A(new_n2177_), .B1(new_n2251_), .B2(new_n2253_), .ZN(new_n2254_));
  NAND2_X1  g2062(.A1(new_n2246_), .A2(new_n2247_), .ZN(new_n2255_));
  NAND2_X1  g2063(.A1(new_n2252_), .A2(new_n2249_), .ZN(new_n2256_));
  NAND2_X1  g2064(.A1(new_n2255_), .A2(new_n2256_), .ZN(new_n2257_));
  NAND3_X1  g2065(.A1(new_n2257_), .A2(new_n2176_), .A3(new_n2250_), .ZN(new_n2258_));
  NOR2_X1   g2066(.A1(new_n310_), .A2(new_n1438_), .ZN(new_n2259_));
  INV_X1    g2067(.A(new_n2259_), .ZN(new_n2260_));
  NAND3_X1  g2068(.A1(new_n2254_), .A2(new_n2258_), .A3(new_n2260_), .ZN(new_n2261_));
  INV_X1    g2069(.A(new_n2261_), .ZN(new_n2262_));
  INV_X1    g2070(.A(new_n2146_), .ZN(new_n2263_));
  NAND2_X1  g2071(.A1(new_n2263_), .A2(new_n2144_), .ZN(new_n2264_));
  INV_X1    g2072(.A(new_n2264_), .ZN(new_n2265_));
  AOI21_X1  g2073(.A(new_n2260_), .B1(new_n2254_), .B2(new_n2258_), .ZN(new_n2266_));
  NOR3_X1   g2074(.A1(new_n2262_), .A2(new_n2265_), .A3(new_n2266_), .ZN(new_n2267_));
  INV_X1    g2075(.A(new_n2266_), .ZN(new_n2268_));
  AOI21_X1  g2076(.A(new_n2264_), .B1(new_n2268_), .B2(new_n2261_), .ZN(new_n2269_));
  OAI21_X1  g2077(.A(new_n2175_), .B1(new_n2267_), .B2(new_n2269_), .ZN(new_n2270_));
  OAI21_X1  g2078(.A(new_n2265_), .B1(new_n2262_), .B2(new_n2266_), .ZN(new_n2271_));
  NAND3_X1  g2079(.A1(new_n2268_), .A2(new_n2261_), .A3(new_n2264_), .ZN(new_n2272_));
  OAI211_X1 g2080(.A(new_n2271_), .B(new_n2272_), .C1(new_n241_), .C2(new_n1654_), .ZN(new_n2273_));
  NAND2_X1  g2081(.A1(new_n2270_), .A2(new_n2273_), .ZN(new_n2274_));
  NAND2_X1  g2082(.A1(new_n2157_), .A2(new_n2151_), .ZN(new_n2275_));
  XNOR2_X1  g2083(.A(new_n2274_), .B(new_n2275_), .ZN(new_n2276_));
  XNOR2_X1  g2084(.A(new_n2174_), .B(new_n2276_), .ZN(G6180gat));
  AOI21_X1  g2085(.A(new_n2274_), .B1(new_n2151_), .B2(new_n2157_), .ZN(new_n2278_));
  AOI21_X1  g2086(.A(new_n2278_), .B1(new_n2174_), .B2(new_n2276_), .ZN(new_n2279_));
  NAND2_X1  g2087(.A1(new_n2234_), .A2(new_n2233_), .ZN(new_n2280_));
  AND2_X1   g2088(.A1(new_n2227_), .A2(new_n2222_), .ZN(new_n2281_));
  INV_X1    g2089(.A(KEYINPUT94), .ZN(new_n2282_));
  AND2_X1   g2090(.A1(new_n2204_), .A2(new_n2202_), .ZN(new_n2283_));
  NAND2_X1  g2091(.A1(new_n2199_), .A2(new_n2200_), .ZN(new_n2284_));
  NAND2_X1  g2092(.A1(new_n2284_), .A2(new_n2196_), .ZN(new_n2285_));
  INV_X1    g2093(.A(new_n2192_), .ZN(new_n2286_));
  NAND2_X1  g2094(.A1(new_n2286_), .A2(new_n2193_), .ZN(new_n2287_));
  NAND2_X1  g2095(.A1(new_n2287_), .A2(KEYINPUT92), .ZN(new_n2288_));
  INV_X1    g2096(.A(KEYINPUT92), .ZN(new_n2289_));
  NAND3_X1  g2097(.A1(new_n2286_), .A2(new_n2289_), .A3(new_n2193_), .ZN(new_n2290_));
  NAND3_X1  g2098(.A1(new_n2288_), .A2(new_n2191_), .A3(new_n2290_), .ZN(new_n2291_));
  OR3_X1    g2099(.A1(new_n2291_), .A2(new_n1872_), .A3(new_n300_), .ZN(new_n2292_));
  NOR2_X1   g2100(.A1(new_n1676_), .A2(new_n355_), .ZN(new_n2293_));
  INV_X1    g2101(.A(new_n2293_), .ZN(new_n2294_));
  OAI21_X1  g2102(.A(new_n2291_), .B1(new_n1872_), .B2(new_n300_), .ZN(new_n2295_));
  NAND3_X1  g2103(.A1(new_n2292_), .A2(new_n2294_), .A3(new_n2295_), .ZN(new_n2296_));
  INV_X1    g2104(.A(new_n2296_), .ZN(new_n2297_));
  INV_X1    g2105(.A(KEYINPUT93), .ZN(new_n2298_));
  AOI21_X1  g2106(.A(new_n2294_), .B1(new_n2292_), .B2(new_n2295_), .ZN(new_n2299_));
  NOR3_X1   g2107(.A1(new_n2297_), .A2(new_n2298_), .A3(new_n2299_), .ZN(new_n2300_));
  NAND2_X1  g2108(.A1(new_n2292_), .A2(new_n2295_), .ZN(new_n2301_));
  NAND2_X1  g2109(.A1(new_n2301_), .A2(new_n2293_), .ZN(new_n2302_));
  AOI21_X1  g2110(.A(KEYINPUT93), .B1(new_n2302_), .B2(new_n2296_), .ZN(new_n2303_));
  OAI21_X1  g2111(.A(new_n2285_), .B1(new_n2300_), .B2(new_n2303_), .ZN(new_n2304_));
  OAI21_X1  g2112(.A(new_n2298_), .B1(new_n2297_), .B2(new_n2299_), .ZN(new_n2305_));
  NAND3_X1  g2113(.A1(new_n2302_), .A2(KEYINPUT93), .A3(new_n2296_), .ZN(new_n2306_));
  NAND4_X1  g2114(.A1(new_n2305_), .A2(new_n2306_), .A3(new_n2196_), .A4(new_n2284_), .ZN(new_n2307_));
  NAND2_X1  g2115(.A1(new_n2304_), .A2(new_n2307_), .ZN(new_n2308_));
  NOR2_X1   g2116(.A1(new_n1681_), .A2(new_n601_), .ZN(new_n2309_));
  NAND2_X1  g2117(.A1(new_n2308_), .A2(new_n2309_), .ZN(new_n2310_));
  OAI211_X1 g2118(.A(new_n2304_), .B(new_n2307_), .C1(new_n1681_), .C2(new_n601_), .ZN(new_n2311_));
  NAND2_X1  g2119(.A1(new_n2310_), .A2(new_n2311_), .ZN(new_n2312_));
  OR2_X1    g2120(.A1(new_n2283_), .A2(new_n2312_), .ZN(new_n2313_));
  NOR2_X1   g2121(.A1(new_n944_), .A2(new_n613_), .ZN(new_n2314_));
  INV_X1    g2122(.A(new_n2314_), .ZN(new_n2315_));
  NAND2_X1  g2123(.A1(new_n2283_), .A2(new_n2312_), .ZN(new_n2316_));
  NAND3_X1  g2124(.A1(new_n2313_), .A2(new_n2315_), .A3(new_n2316_), .ZN(new_n2317_));
  INV_X1    g2125(.A(new_n2317_), .ZN(new_n2318_));
  AOI21_X1  g2126(.A(new_n2315_), .B1(new_n2313_), .B2(new_n2316_), .ZN(new_n2319_));
  OAI21_X1  g2127(.A(new_n2282_), .B1(new_n2318_), .B2(new_n2319_), .ZN(new_n2320_));
  INV_X1    g2128(.A(new_n2319_), .ZN(new_n2321_));
  NAND3_X1  g2129(.A1(new_n2321_), .A2(KEYINPUT94), .A3(new_n2317_), .ZN(new_n2322_));
  INV_X1    g2130(.A(new_n2207_), .ZN(new_n2323_));
  NAND2_X1  g2131(.A1(new_n2210_), .A2(new_n2323_), .ZN(new_n2324_));
  NAND3_X1  g2132(.A1(new_n2320_), .A2(new_n2322_), .A3(new_n2324_), .ZN(new_n2325_));
  NAND2_X1  g2133(.A1(new_n2321_), .A2(new_n2317_), .ZN(new_n2326_));
  NAND4_X1  g2134(.A1(new_n2326_), .A2(new_n2282_), .A3(new_n2323_), .A4(new_n2210_), .ZN(new_n2327_));
  NAND2_X1  g2135(.A1(G188gat), .A2(G426gat), .ZN(new_n2328_));
  NAND3_X1  g2136(.A1(new_n2325_), .A2(new_n2327_), .A3(new_n2328_), .ZN(new_n2329_));
  INV_X1    g2137(.A(new_n2329_), .ZN(new_n2330_));
  AOI21_X1  g2138(.A(new_n2328_), .B1(new_n2325_), .B2(new_n2327_), .ZN(new_n2331_));
  NOR2_X1   g2139(.A1(new_n2330_), .A2(new_n2331_), .ZN(new_n2332_));
  NOR2_X1   g2140(.A1(new_n2218_), .A2(new_n2215_), .ZN(new_n2333_));
  INV_X1    g2141(.A(new_n2333_), .ZN(new_n2334_));
  NAND2_X1  g2142(.A1(new_n2332_), .A2(new_n2334_), .ZN(new_n2335_));
  OAI21_X1  g2143(.A(new_n2333_), .B1(new_n2330_), .B2(new_n2331_), .ZN(new_n2336_));
  NAND2_X1  g2144(.A1(new_n2335_), .A2(new_n2336_), .ZN(new_n2337_));
  NOR2_X1   g2145(.A1(new_n799_), .A2(new_n768_), .ZN(new_n2338_));
  NOR2_X1   g2146(.A1(new_n2337_), .A2(new_n2338_), .ZN(new_n2339_));
  AND2_X1   g2147(.A1(new_n2337_), .A2(new_n2338_), .ZN(new_n2340_));
  OR3_X1    g2148(.A1(new_n2281_), .A2(new_n2339_), .A3(new_n2340_), .ZN(new_n2341_));
  OAI21_X1  g2149(.A(new_n2281_), .B1(new_n2339_), .B2(new_n2340_), .ZN(new_n2342_));
  NAND2_X1  g2150(.A1(G154gat), .A2(G460gat), .ZN(new_n2343_));
  NAND2_X1  g2151(.A1(new_n2343_), .A2(KEYINPUT95), .ZN(new_n2344_));
  NAND3_X1  g2152(.A1(new_n2341_), .A2(new_n2342_), .A3(new_n2344_), .ZN(new_n2345_));
  INV_X1    g2153(.A(new_n2345_), .ZN(new_n2346_));
  OR2_X1    g2154(.A1(new_n2343_), .A2(KEYINPUT95), .ZN(new_n2347_));
  AOI22_X1  g2155(.A1(new_n2341_), .A2(new_n2342_), .B1(new_n2344_), .B2(new_n2347_), .ZN(new_n2348_));
  OAI21_X1  g2156(.A(new_n2280_), .B1(new_n2346_), .B2(new_n2348_), .ZN(new_n2349_));
  NAND2_X1  g2157(.A1(new_n2341_), .A2(new_n2342_), .ZN(new_n2350_));
  NAND2_X1  g2158(.A1(new_n2347_), .A2(new_n2344_), .ZN(new_n2351_));
  NAND2_X1  g2159(.A1(new_n2350_), .A2(new_n2351_), .ZN(new_n2352_));
  NAND4_X1  g2160(.A1(new_n2352_), .A2(new_n2233_), .A3(new_n2234_), .A4(new_n2345_), .ZN(new_n2353_));
  NAND2_X1  g2161(.A1(new_n2349_), .A2(new_n2353_), .ZN(new_n2354_));
  NOR2_X1   g2162(.A1(new_n651_), .A2(new_n1419_), .ZN(new_n2355_));
  NAND2_X1  g2163(.A1(new_n2354_), .A2(new_n2355_), .ZN(new_n2356_));
  XOR2_X1   g2164(.A(new_n2355_), .B(KEYINPUT96), .Z(new_n2357_));
  NAND3_X1  g2165(.A1(new_n2349_), .A2(new_n2353_), .A3(new_n2357_), .ZN(new_n2358_));
  NAND2_X1  g2166(.A1(new_n2356_), .A2(new_n2358_), .ZN(new_n2359_));
  NAND3_X1  g2167(.A1(new_n2237_), .A2(G120gat), .A3(G477gat), .ZN(new_n2360_));
  NAND2_X1  g2168(.A1(new_n2360_), .A2(new_n2238_), .ZN(new_n2361_));
  NAND2_X1  g2169(.A1(new_n2359_), .A2(new_n2361_), .ZN(new_n2362_));
  NAND2_X1  g2170(.A1(G120gat), .A2(G494gat), .ZN(new_n2363_));
  NAND4_X1  g2171(.A1(new_n2356_), .A2(new_n2238_), .A3(new_n2358_), .A4(new_n2360_), .ZN(new_n2364_));
  NAND3_X1  g2172(.A1(new_n2362_), .A2(new_n2363_), .A3(new_n2364_), .ZN(new_n2365_));
  INV_X1    g2173(.A(new_n2365_), .ZN(new_n2366_));
  AOI21_X1  g2174(.A(new_n2363_), .B1(new_n2362_), .B2(new_n2364_), .ZN(new_n2367_));
  NOR2_X1   g2175(.A1(new_n2366_), .A2(new_n2367_), .ZN(new_n2368_));
  NAND2_X1  g2176(.A1(new_n2247_), .A2(new_n2248_), .ZN(new_n2369_));
  NAND2_X1  g2177(.A1(new_n2369_), .A2(new_n2246_), .ZN(new_n2370_));
  OR2_X1    g2178(.A1(new_n2368_), .A2(new_n2370_), .ZN(new_n2371_));
  NAND2_X1  g2179(.A1(new_n2368_), .A2(new_n2370_), .ZN(new_n2372_));
  NAND2_X1  g2180(.A1(new_n2371_), .A2(new_n2372_), .ZN(new_n2373_));
  NAND3_X1  g2181(.A1(new_n2373_), .A2(G103gat), .A3(G511gat), .ZN(new_n2374_));
  NAND2_X1  g2182(.A1(G103gat), .A2(G511gat), .ZN(new_n2375_));
  NAND3_X1  g2183(.A1(new_n2371_), .A2(new_n2375_), .A3(new_n2372_), .ZN(new_n2376_));
  NAND2_X1  g2184(.A1(new_n2374_), .A2(new_n2376_), .ZN(new_n2377_));
  NAND3_X1  g2185(.A1(new_n2377_), .A2(new_n2254_), .A3(new_n2261_), .ZN(new_n2378_));
  NAND2_X1  g2186(.A1(G86gat), .A2(G528gat), .ZN(new_n2379_));
  NAND2_X1  g2187(.A1(new_n2261_), .A2(new_n2254_), .ZN(new_n2380_));
  NAND3_X1  g2188(.A1(new_n2374_), .A2(new_n2380_), .A3(new_n2376_), .ZN(new_n2381_));
  NAND3_X1  g2189(.A1(new_n2378_), .A2(new_n2379_), .A3(new_n2381_), .ZN(new_n2382_));
  INV_X1    g2190(.A(new_n2382_), .ZN(new_n2383_));
  AOI21_X1  g2191(.A(new_n2379_), .B1(new_n2378_), .B2(new_n2381_), .ZN(new_n2384_));
  OAI211_X1 g2192(.A(new_n2272_), .B(new_n2273_), .C1(new_n2383_), .C2(new_n2384_), .ZN(new_n2385_));
  INV_X1    g2193(.A(new_n2384_), .ZN(new_n2386_));
  NAND2_X1  g2194(.A1(new_n2273_), .A2(new_n2272_), .ZN(new_n2387_));
  NAND3_X1  g2195(.A1(new_n2386_), .A2(new_n2387_), .A3(new_n2382_), .ZN(new_n2388_));
  NAND2_X1  g2196(.A1(new_n2385_), .A2(new_n2388_), .ZN(new_n2389_));
  XNOR2_X1  g2197(.A(new_n2279_), .B(new_n2389_), .ZN(G6190gat));
  OAI21_X1  g2198(.A(new_n2388_), .B1(new_n2279_), .B2(new_n2389_), .ZN(new_n2391_));
  XNOR2_X1  g2199(.A(new_n2391_), .B(KEYINPUT106), .ZN(new_n2392_));
  NOR2_X1   g2200(.A1(new_n452_), .A2(new_n1654_), .ZN(new_n2393_));
  INV_X1    g2201(.A(new_n2364_), .ZN(new_n2394_));
  AOI21_X1  g2202(.A(new_n2394_), .B1(new_n2363_), .B2(new_n2362_), .ZN(new_n2395_));
  INV_X1    g2203(.A(new_n2395_), .ZN(new_n2396_));
  INV_X1    g2204(.A(KEYINPUT101), .ZN(new_n2397_));
  NOR2_X1   g2205(.A1(new_n799_), .A2(new_n918_), .ZN(new_n2398_));
  NAND3_X1  g2206(.A1(new_n2324_), .A2(new_n2317_), .A3(new_n2321_), .ZN(new_n2399_));
  NAND2_X1  g2207(.A1(new_n2329_), .A2(new_n2399_), .ZN(new_n2400_));
  NOR3_X1   g2208(.A1(new_n2300_), .A2(new_n2303_), .A3(new_n2285_), .ZN(new_n2401_));
  OAI21_X1  g2209(.A(new_n2304_), .B1(new_n2401_), .B2(new_n2309_), .ZN(new_n2402_));
  INV_X1    g2210(.A(KEYINPUT98), .ZN(new_n2403_));
  NAND2_X1  g2211(.A1(new_n2402_), .A2(new_n2403_), .ZN(new_n2404_));
  OAI211_X1 g2212(.A(KEYINPUT98), .B(new_n2304_), .C1(new_n2401_), .C2(new_n2309_), .ZN(new_n2405_));
  NAND2_X1  g2213(.A1(new_n2404_), .A2(new_n2405_), .ZN(new_n2406_));
  NAND2_X1  g2214(.A1(new_n2296_), .A2(new_n2295_), .ZN(new_n2407_));
  NOR2_X1   g2215(.A1(new_n1872_), .A2(new_n355_), .ZN(new_n2408_));
  NAND2_X1  g2216(.A1(new_n2407_), .A2(new_n2408_), .ZN(new_n2409_));
  XOR2_X1   g2217(.A(new_n2408_), .B(KEYINPUT97), .Z(new_n2410_));
  OAI21_X1  g2218(.A(new_n2409_), .B1(new_n2407_), .B2(new_n2410_), .ZN(new_n2411_));
  NOR2_X1   g2219(.A1(new_n1676_), .A2(new_n601_), .ZN(new_n2412_));
  XNOR2_X1  g2220(.A(new_n2411_), .B(new_n2412_), .ZN(new_n2413_));
  NAND2_X1  g2221(.A1(new_n2406_), .A2(new_n2413_), .ZN(new_n2414_));
  NAND2_X1  g2222(.A1(G222gat), .A2(G409gat), .ZN(new_n2415_));
  INV_X1    g2223(.A(new_n2413_), .ZN(new_n2416_));
  NAND3_X1  g2224(.A1(new_n2404_), .A2(new_n2416_), .A3(new_n2405_), .ZN(new_n2417_));
  NAND3_X1  g2225(.A1(new_n2414_), .A2(new_n2415_), .A3(new_n2417_), .ZN(new_n2418_));
  INV_X1    g2226(.A(new_n2418_), .ZN(new_n2419_));
  AOI21_X1  g2227(.A(new_n2415_), .B1(new_n2414_), .B2(new_n2417_), .ZN(new_n2420_));
  NOR2_X1   g2228(.A1(new_n2419_), .A2(new_n2420_), .ZN(new_n2421_));
  NAND2_X1  g2229(.A1(new_n2317_), .A2(new_n2313_), .ZN(new_n2422_));
  NAND2_X1  g2230(.A1(new_n2421_), .A2(new_n2422_), .ZN(new_n2423_));
  OAI211_X1 g2231(.A(new_n2313_), .B(new_n2317_), .C1(new_n2419_), .C2(new_n2420_), .ZN(new_n2424_));
  OAI211_X1 g2232(.A(new_n2423_), .B(new_n2424_), .C1(new_n944_), .C2(new_n624_), .ZN(new_n2425_));
  NAND2_X1  g2233(.A1(new_n2423_), .A2(new_n2424_), .ZN(new_n2426_));
  NOR2_X1   g2234(.A1(new_n944_), .A2(new_n624_), .ZN(new_n2427_));
  NAND2_X1  g2235(.A1(new_n2426_), .A2(new_n2427_), .ZN(new_n2428_));
  NAND3_X1  g2236(.A1(new_n2400_), .A2(new_n2425_), .A3(new_n2428_), .ZN(new_n2429_));
  NAND2_X1  g2237(.A1(new_n2428_), .A2(new_n2425_), .ZN(new_n2430_));
  NAND3_X1  g2238(.A1(new_n2430_), .A2(new_n2329_), .A3(new_n2399_), .ZN(new_n2431_));
  NAND2_X1  g2239(.A1(new_n2429_), .A2(new_n2431_), .ZN(new_n2432_));
  NOR2_X1   g2240(.A1(new_n1093_), .A2(new_n768_), .ZN(new_n2433_));
  NAND2_X1  g2241(.A1(new_n2432_), .A2(new_n2433_), .ZN(new_n2434_));
  OAI211_X1 g2242(.A(new_n2429_), .B(new_n2431_), .C1(new_n1093_), .C2(new_n768_), .ZN(new_n2435_));
  NAND2_X1  g2243(.A1(new_n2434_), .A2(new_n2435_), .ZN(new_n2436_));
  INV_X1    g2244(.A(new_n2336_), .ZN(new_n2437_));
  OAI211_X1 g2245(.A(KEYINPUT99), .B(new_n2335_), .C1(new_n2437_), .C2(new_n2338_), .ZN(new_n2438_));
  NAND2_X1  g2246(.A1(new_n2436_), .A2(new_n2438_), .ZN(new_n2439_));
  OAI21_X1  g2247(.A(new_n2335_), .B1(new_n2437_), .B2(new_n2338_), .ZN(new_n2440_));
  INV_X1    g2248(.A(KEYINPUT99), .ZN(new_n2441_));
  NAND2_X1  g2249(.A1(new_n2440_), .A2(new_n2441_), .ZN(new_n2442_));
  AND2_X1   g2250(.A1(new_n2442_), .A2(new_n2438_), .ZN(new_n2443_));
  OAI211_X1 g2251(.A(new_n2398_), .B(new_n2439_), .C1(new_n2443_), .C2(new_n2436_), .ZN(new_n2444_));
  INV_X1    g2252(.A(new_n2398_), .ZN(new_n2445_));
  AOI21_X1  g2253(.A(new_n2436_), .B1(new_n2442_), .B2(new_n2438_), .ZN(new_n2446_));
  AND2_X1   g2254(.A1(new_n2436_), .A2(new_n2438_), .ZN(new_n2447_));
  OAI21_X1  g2255(.A(new_n2445_), .B1(new_n2446_), .B2(new_n2447_), .ZN(new_n2448_));
  NAND3_X1  g2256(.A1(new_n2444_), .A2(KEYINPUT100), .A3(new_n2448_), .ZN(new_n2449_));
  INV_X1    g2257(.A(new_n2449_), .ZN(new_n2450_));
  AOI21_X1  g2258(.A(KEYINPUT100), .B1(new_n2444_), .B2(new_n2448_), .ZN(new_n2451_));
  OAI21_X1  g2259(.A(new_n2397_), .B1(new_n2450_), .B2(new_n2451_), .ZN(new_n2452_));
  INV_X1    g2260(.A(new_n2451_), .ZN(new_n2453_));
  NAND3_X1  g2261(.A1(new_n2453_), .A2(KEYINPUT101), .A3(new_n2449_), .ZN(new_n2454_));
  NAND2_X1  g2262(.A1(new_n2452_), .A2(new_n2454_), .ZN(new_n2455_));
  NAND3_X1  g2263(.A1(new_n2341_), .A2(G154gat), .A3(G460gat), .ZN(new_n2456_));
  NAND2_X1  g2264(.A1(new_n2456_), .A2(new_n2342_), .ZN(new_n2457_));
  INV_X1    g2265(.A(new_n2457_), .ZN(new_n2458_));
  NAND2_X1  g2266(.A1(new_n2455_), .A2(new_n2458_), .ZN(new_n2459_));
  NOR2_X1   g2267(.A1(new_n960_), .A2(new_n1419_), .ZN(new_n2460_));
  NAND2_X1  g2268(.A1(new_n2452_), .A2(new_n2457_), .ZN(new_n2461_));
  NAND3_X1  g2269(.A1(new_n2459_), .A2(new_n2460_), .A3(new_n2461_), .ZN(new_n2462_));
  INV_X1    g2270(.A(new_n2460_), .ZN(new_n2463_));
  AOI21_X1  g2271(.A(new_n2457_), .B1(new_n2452_), .B2(new_n2454_), .ZN(new_n2464_));
  NAND2_X1  g2272(.A1(new_n2453_), .A2(new_n2449_), .ZN(new_n2465_));
  AOI21_X1  g2273(.A(new_n2458_), .B1(new_n2465_), .B2(new_n2397_), .ZN(new_n2466_));
  OAI21_X1  g2274(.A(new_n2463_), .B1(new_n2464_), .B2(new_n2466_), .ZN(new_n2467_));
  NAND2_X1  g2275(.A1(new_n2358_), .A2(new_n2349_), .ZN(new_n2468_));
  AND3_X1   g2276(.A1(new_n2462_), .A2(new_n2467_), .A3(new_n2468_), .ZN(new_n2469_));
  AOI21_X1  g2277(.A(new_n2468_), .B1(new_n2462_), .B2(new_n2467_), .ZN(new_n2470_));
  NOR2_X1   g2278(.A1(new_n651_), .A2(new_n1426_), .ZN(new_n2471_));
  NOR3_X1   g2279(.A1(new_n2469_), .A2(new_n2470_), .A3(new_n2471_), .ZN(new_n2472_));
  INV_X1    g2280(.A(new_n2471_), .ZN(new_n2473_));
  INV_X1    g2281(.A(new_n2468_), .ZN(new_n2474_));
  AOI21_X1  g2282(.A(new_n2460_), .B1(new_n2459_), .B2(new_n2461_), .ZN(new_n2475_));
  NOR3_X1   g2283(.A1(new_n2464_), .A2(new_n2466_), .A3(new_n2463_), .ZN(new_n2476_));
  OAI21_X1  g2284(.A(new_n2474_), .B1(new_n2475_), .B2(new_n2476_), .ZN(new_n2477_));
  NAND3_X1  g2285(.A1(new_n2462_), .A2(new_n2467_), .A3(new_n2468_), .ZN(new_n2478_));
  AOI21_X1  g2286(.A(new_n2473_), .B1(new_n2477_), .B2(new_n2478_), .ZN(new_n2479_));
  OAI21_X1  g2287(.A(new_n2396_), .B1(new_n2472_), .B2(new_n2479_), .ZN(new_n2480_));
  INV_X1    g2288(.A(KEYINPUT103), .ZN(new_n2481_));
  NAND2_X1  g2289(.A1(new_n2480_), .A2(new_n2481_), .ZN(new_n2482_));
  OAI21_X1  g2290(.A(new_n2471_), .B1(new_n2469_), .B2(new_n2470_), .ZN(new_n2483_));
  NAND3_X1  g2291(.A1(new_n2477_), .A2(new_n2473_), .A3(new_n2478_), .ZN(new_n2484_));
  NAND2_X1  g2292(.A1(new_n2483_), .A2(new_n2484_), .ZN(new_n2485_));
  NAND3_X1  g2293(.A1(new_n2485_), .A2(KEYINPUT103), .A3(new_n2396_), .ZN(new_n2486_));
  NAND2_X1  g2294(.A1(new_n2482_), .A2(new_n2486_), .ZN(new_n2487_));
  NOR2_X1   g2295(.A1(new_n532_), .A2(new_n1438_), .ZN(new_n2488_));
  NAND3_X1  g2296(.A1(new_n2483_), .A2(new_n2395_), .A3(new_n2484_), .ZN(new_n2489_));
  NAND2_X1  g2297(.A1(new_n2489_), .A2(KEYINPUT102), .ZN(new_n2490_));
  INV_X1    g2298(.A(KEYINPUT102), .ZN(new_n2491_));
  NAND4_X1  g2299(.A1(new_n2483_), .A2(new_n2484_), .A3(new_n2491_), .A4(new_n2395_), .ZN(new_n2492_));
  NAND2_X1  g2300(.A1(new_n2490_), .A2(new_n2492_), .ZN(new_n2493_));
  AND3_X1   g2301(.A1(new_n2487_), .A2(new_n2488_), .A3(new_n2493_), .ZN(new_n2494_));
  AOI21_X1  g2302(.A(new_n2488_), .B1(new_n2487_), .B2(new_n2493_), .ZN(new_n2495_));
  NAND2_X1  g2303(.A1(new_n2376_), .A2(new_n2372_), .ZN(new_n2496_));
  INV_X1    g2304(.A(new_n2496_), .ZN(new_n2497_));
  NOR3_X1   g2305(.A1(new_n2494_), .A2(new_n2495_), .A3(new_n2497_), .ZN(new_n2498_));
  AND2_X1   g2306(.A1(new_n2489_), .A2(KEYINPUT102), .ZN(new_n2499_));
  INV_X1    g2307(.A(new_n2492_), .ZN(new_n2500_));
  AOI21_X1  g2308(.A(KEYINPUT103), .B1(new_n2485_), .B2(new_n2396_), .ZN(new_n2501_));
  AOI211_X1 g2309(.A(new_n2481_), .B(new_n2395_), .C1(new_n2483_), .C2(new_n2484_), .ZN(new_n2502_));
  OAI22_X1  g2310(.A1(new_n2499_), .A2(new_n2500_), .B1(new_n2501_), .B2(new_n2502_), .ZN(new_n2503_));
  INV_X1    g2311(.A(new_n2488_), .ZN(new_n2504_));
  NAND2_X1  g2312(.A1(new_n2503_), .A2(new_n2504_), .ZN(new_n2505_));
  NAND3_X1  g2313(.A1(new_n2487_), .A2(new_n2488_), .A3(new_n2493_), .ZN(new_n2506_));
  AOI21_X1  g2314(.A(new_n2496_), .B1(new_n2505_), .B2(new_n2506_), .ZN(new_n2507_));
  OAI21_X1  g2315(.A(new_n2393_), .B1(new_n2498_), .B2(new_n2507_), .ZN(new_n2508_));
  OAI21_X1  g2316(.A(new_n2497_), .B1(new_n2494_), .B2(new_n2495_), .ZN(new_n2509_));
  NAND3_X1  g2317(.A1(new_n2505_), .A2(new_n2496_), .A3(new_n2506_), .ZN(new_n2510_));
  INV_X1    g2318(.A(new_n2393_), .ZN(new_n2511_));
  NAND3_X1  g2319(.A1(new_n2509_), .A2(new_n2510_), .A3(new_n2511_), .ZN(new_n2512_));
  INV_X1    g2320(.A(new_n2381_), .ZN(new_n2513_));
  AOI21_X1  g2321(.A(new_n2513_), .B1(new_n2378_), .B2(new_n2379_), .ZN(new_n2514_));
  NAND3_X1  g2322(.A1(new_n2508_), .A2(new_n2512_), .A3(new_n2514_), .ZN(new_n2515_));
  INV_X1    g2323(.A(KEYINPUT105), .ZN(new_n2516_));
  NAND2_X1  g2324(.A1(new_n2515_), .A2(new_n2516_), .ZN(new_n2517_));
  NAND4_X1  g2325(.A1(new_n2508_), .A2(KEYINPUT105), .A3(new_n2512_), .A4(new_n2514_), .ZN(new_n2518_));
  NAND2_X1  g2326(.A1(new_n2517_), .A2(new_n2518_), .ZN(new_n2519_));
  NAND2_X1  g2327(.A1(new_n2509_), .A2(new_n2510_), .ZN(new_n2520_));
  AOI21_X1  g2328(.A(new_n2514_), .B1(KEYINPUT104), .B2(new_n2520_), .ZN(new_n2521_));
  NAND2_X1  g2329(.A1(new_n2508_), .A2(new_n2512_), .ZN(new_n2522_));
  OAI21_X1  g2330(.A(new_n2521_), .B1(new_n2522_), .B2(KEYINPUT104), .ZN(new_n2523_));
  NAND2_X1  g2331(.A1(new_n2519_), .A2(new_n2523_), .ZN(new_n2524_));
  XNOR2_X1  g2332(.A(new_n2392_), .B(new_n2524_), .ZN(G6200gat));
  NOR2_X1   g2333(.A1(new_n2522_), .A2(new_n2514_), .ZN(new_n2526_));
  AOI21_X1  g2334(.A(new_n2526_), .B1(new_n2391_), .B2(new_n2524_), .ZN(new_n2527_));
  NAND2_X1  g2335(.A1(new_n2512_), .A2(new_n2510_), .ZN(new_n2528_));
  INV_X1    g2336(.A(new_n2528_), .ZN(new_n2529_));
  NOR2_X1   g2337(.A1(new_n651_), .A2(new_n1438_), .ZN(new_n2530_));
  INV_X1    g2338(.A(KEYINPUT109), .ZN(new_n2531_));
  AOI22_X1  g2339(.A1(new_n2418_), .A2(KEYINPUT107), .B1(new_n2406_), .B2(new_n2413_), .ZN(new_n2532_));
  OAI21_X1  g2340(.A(new_n2532_), .B1(KEYINPUT107), .B2(new_n2418_), .ZN(new_n2533_));
  OAI21_X1  g2341(.A(new_n2411_), .B1(new_n1676_), .B2(new_n601_), .ZN(new_n2534_));
  AND2_X1   g2342(.A1(new_n2296_), .A2(new_n2295_), .ZN(new_n2535_));
  OAI21_X1  g2343(.A(new_n2534_), .B1(new_n2535_), .B2(new_n2410_), .ZN(new_n2536_));
  NAND2_X1  g2344(.A1(G256gat), .A2(G392gat), .ZN(new_n2537_));
  XNOR2_X1  g2345(.A(new_n2536_), .B(new_n2537_), .ZN(new_n2538_));
  NOR2_X1   g2346(.A1(new_n1676_), .A2(new_n613_), .ZN(new_n2539_));
  OR2_X1    g2347(.A1(new_n2538_), .A2(new_n2539_), .ZN(new_n2540_));
  NAND2_X1  g2348(.A1(new_n2538_), .A2(new_n2539_), .ZN(new_n2541_));
  NAND3_X1  g2349(.A1(new_n2533_), .A2(new_n2540_), .A3(new_n2541_), .ZN(new_n2542_));
  NAND2_X1  g2350(.A1(new_n2540_), .A2(new_n2541_), .ZN(new_n2543_));
  NAND3_X1  g2351(.A1(new_n2543_), .A2(new_n2414_), .A3(new_n2418_), .ZN(new_n2544_));
  NAND2_X1  g2352(.A1(new_n2542_), .A2(new_n2544_), .ZN(new_n2545_));
  NAND3_X1  g2353(.A1(new_n2545_), .A2(G222gat), .A3(G426gat), .ZN(new_n2546_));
  OAI211_X1 g2354(.A(new_n2542_), .B(new_n2544_), .C1(new_n1681_), .C2(new_n624_), .ZN(new_n2547_));
  NAND2_X1  g2355(.A1(new_n2546_), .A2(new_n2547_), .ZN(new_n2548_));
  AND2_X1   g2356(.A1(new_n2425_), .A2(new_n2423_), .ZN(new_n2549_));
  OR2_X1    g2357(.A1(new_n2548_), .A2(new_n2549_), .ZN(new_n2550_));
  NAND2_X1  g2358(.A1(new_n2548_), .A2(new_n2549_), .ZN(new_n2551_));
  NAND2_X1  g2359(.A1(new_n2550_), .A2(new_n2551_), .ZN(new_n2552_));
  INV_X1    g2360(.A(new_n2552_), .ZN(new_n2553_));
  NAND2_X1  g2361(.A1(G205gat), .A2(G443gat), .ZN(new_n2554_));
  INV_X1    g2362(.A(KEYINPUT108), .ZN(new_n2555_));
  NOR2_X1   g2363(.A1(new_n2554_), .A2(new_n2555_), .ZN(new_n2556_));
  NOR2_X1   g2364(.A1(new_n2553_), .A2(new_n2556_), .ZN(new_n2557_));
  INV_X1    g2365(.A(new_n2556_), .ZN(new_n2558_));
  NAND2_X1  g2366(.A1(new_n2554_), .A2(new_n2555_), .ZN(new_n2559_));
  AOI21_X1  g2367(.A(new_n2552_), .B1(new_n2558_), .B2(new_n2559_), .ZN(new_n2560_));
  OAI21_X1  g2368(.A(new_n2531_), .B1(new_n2557_), .B2(new_n2560_), .ZN(new_n2561_));
  NAND2_X1  g2369(.A1(new_n2558_), .A2(new_n2559_), .ZN(new_n2562_));
  NAND2_X1  g2370(.A1(new_n2553_), .A2(new_n2562_), .ZN(new_n2563_));
  OAI211_X1 g2371(.A(new_n2563_), .B(KEYINPUT109), .C1(new_n2553_), .C2(new_n2556_), .ZN(new_n2564_));
  NAND2_X1  g2372(.A1(new_n2561_), .A2(new_n2564_), .ZN(new_n2565_));
  AND2_X1   g2373(.A1(new_n2435_), .A2(new_n2429_), .ZN(new_n2566_));
  OR2_X1    g2374(.A1(new_n2565_), .A2(new_n2566_), .ZN(new_n2567_));
  NOR2_X1   g2375(.A1(new_n1093_), .A2(new_n918_), .ZN(new_n2568_));
  INV_X1    g2376(.A(new_n2568_), .ZN(new_n2569_));
  OAI211_X1 g2377(.A(new_n2563_), .B(new_n2566_), .C1(new_n2553_), .C2(new_n2556_), .ZN(new_n2570_));
  NAND3_X1  g2378(.A1(new_n2567_), .A2(new_n2569_), .A3(new_n2570_), .ZN(new_n2571_));
  OAI21_X1  g2379(.A(new_n2570_), .B1(new_n2565_), .B2(new_n2566_), .ZN(new_n2572_));
  NAND2_X1  g2380(.A1(new_n2572_), .A2(new_n2568_), .ZN(new_n2573_));
  AND3_X1   g2381(.A1(new_n2571_), .A2(KEYINPUT110), .A3(new_n2573_), .ZN(new_n2574_));
  AOI21_X1  g2382(.A(KEYINPUT110), .B1(new_n2571_), .B2(new_n2573_), .ZN(new_n2575_));
  NOR2_X1   g2383(.A1(new_n2574_), .A2(new_n2575_), .ZN(new_n2576_));
  NAND3_X1  g2384(.A1(new_n2440_), .A2(new_n2435_), .A3(new_n2434_), .ZN(new_n2577_));
  NAND2_X1  g2385(.A1(new_n2448_), .A2(new_n2577_), .ZN(new_n2578_));
  NOR2_X1   g2386(.A1(new_n799_), .A2(new_n1419_), .ZN(new_n2579_));
  XOR2_X1   g2387(.A(new_n2578_), .B(new_n2579_), .Z(new_n2580_));
  NAND2_X1  g2388(.A1(new_n2576_), .A2(new_n2580_), .ZN(new_n2581_));
  NAND2_X1  g2389(.A1(new_n2571_), .A2(new_n2573_), .ZN(new_n2582_));
  OAI21_X1  g2390(.A(new_n2581_), .B1(new_n2582_), .B2(new_n2580_), .ZN(new_n2583_));
  INV_X1    g2391(.A(new_n2465_), .ZN(new_n2584_));
  AOI21_X1  g2392(.A(new_n2475_), .B1(new_n2458_), .B2(new_n2584_), .ZN(new_n2585_));
  AND2_X1   g2393(.A1(new_n2583_), .A2(new_n2585_), .ZN(new_n2586_));
  NOR2_X1   g2394(.A1(new_n2583_), .A2(new_n2585_), .ZN(new_n2587_));
  NOR2_X1   g2395(.A1(new_n960_), .A2(new_n1426_), .ZN(new_n2588_));
  OR3_X1    g2396(.A1(new_n2586_), .A2(new_n2587_), .A3(new_n2588_), .ZN(new_n2589_));
  OAI21_X1  g2397(.A(new_n2588_), .B1(new_n2586_), .B2(new_n2587_), .ZN(new_n2590_));
  NAND2_X1  g2398(.A1(new_n2589_), .A2(new_n2590_), .ZN(new_n2591_));
  NAND2_X1  g2399(.A1(new_n2484_), .A2(new_n2478_), .ZN(new_n2592_));
  OAI21_X1  g2400(.A(new_n2591_), .B1(KEYINPUT111), .B2(new_n2592_), .ZN(new_n2593_));
  XNOR2_X1  g2401(.A(new_n2592_), .B(KEYINPUT111), .ZN(new_n2594_));
  NAND3_X1  g2402(.A1(new_n2594_), .A2(new_n2589_), .A3(new_n2590_), .ZN(new_n2595_));
  AOI21_X1  g2403(.A(new_n2530_), .B1(new_n2593_), .B2(new_n2595_), .ZN(new_n2596_));
  INV_X1    g2404(.A(new_n2596_), .ZN(new_n2597_));
  NAND3_X1  g2405(.A1(new_n2593_), .A2(new_n2530_), .A3(new_n2595_), .ZN(new_n2598_));
  NAND2_X1  g2406(.A1(new_n2597_), .A2(new_n2598_), .ZN(new_n2599_));
  NAND3_X1  g2407(.A1(new_n2483_), .A2(new_n2396_), .A3(new_n2484_), .ZN(new_n2600_));
  NAND3_X1  g2408(.A1(new_n2599_), .A2(new_n2505_), .A3(new_n2600_), .ZN(new_n2601_));
  NOR2_X1   g2409(.A1(new_n532_), .A2(new_n1654_), .ZN(new_n2602_));
  INV_X1    g2410(.A(new_n2602_), .ZN(new_n2603_));
  NAND2_X1  g2411(.A1(new_n2505_), .A2(new_n2600_), .ZN(new_n2604_));
  NAND3_X1  g2412(.A1(new_n2597_), .A2(new_n2604_), .A3(new_n2598_), .ZN(new_n2605_));
  NAND3_X1  g2413(.A1(new_n2601_), .A2(new_n2603_), .A3(new_n2605_), .ZN(new_n2606_));
  INV_X1    g2414(.A(new_n2606_), .ZN(new_n2607_));
  AOI21_X1  g2415(.A(new_n2603_), .B1(new_n2601_), .B2(new_n2605_), .ZN(new_n2608_));
  OAI21_X1  g2416(.A(new_n2529_), .B1(new_n2607_), .B2(new_n2608_), .ZN(new_n2609_));
  INV_X1    g2417(.A(new_n2608_), .ZN(new_n2610_));
  NAND3_X1  g2418(.A1(new_n2610_), .A2(new_n2528_), .A3(new_n2606_), .ZN(new_n2611_));
  NAND2_X1  g2419(.A1(new_n2609_), .A2(new_n2611_), .ZN(new_n2612_));
  XNOR2_X1  g2420(.A(new_n2527_), .B(new_n2612_), .ZN(G6210gat));
  OAI21_X1  g2421(.A(new_n2611_), .B1(new_n2527_), .B2(new_n2612_), .ZN(new_n2614_));
  OAI21_X1  g2422(.A(new_n2536_), .B1(new_n1872_), .B2(new_n601_), .ZN(new_n2615_));
  NAND2_X1  g2423(.A1(new_n2540_), .A2(new_n2615_), .ZN(new_n2616_));
  OAI21_X1  g2424(.A(new_n2616_), .B1(new_n1872_), .B2(new_n613_), .ZN(new_n2617_));
  NAND4_X1  g2425(.A1(new_n2540_), .A2(G256gat), .A3(G409gat), .A4(new_n2615_), .ZN(new_n2618_));
  NAND2_X1  g2426(.A1(new_n2617_), .A2(new_n2618_), .ZN(new_n2619_));
  NOR2_X1   g2427(.A1(new_n1676_), .A2(new_n624_), .ZN(new_n2620_));
  XNOR2_X1  g2428(.A(new_n2619_), .B(new_n2620_), .ZN(new_n2621_));
  XNOR2_X1  g2429(.A(new_n2621_), .B(KEYINPUT113), .ZN(new_n2622_));
  INV_X1    g2430(.A(KEYINPUT113), .ZN(new_n2623_));
  NOR2_X1   g2431(.A1(new_n2621_), .A2(new_n2623_), .ZN(new_n2624_));
  XNOR2_X1  g2432(.A(new_n2542_), .B(KEYINPUT112), .ZN(new_n2625_));
  NAND2_X1  g2433(.A1(new_n2625_), .A2(new_n2547_), .ZN(new_n2626_));
  MUX2_X1   g2434(.A(new_n2622_), .B(new_n2624_), .S(new_n2626_), .Z(new_n2627_));
  NOR2_X1   g2435(.A1(new_n1681_), .A2(new_n768_), .ZN(new_n2628_));
  XNOR2_X1  g2436(.A(new_n2627_), .B(new_n2628_), .ZN(new_n2629_));
  NOR2_X1   g2437(.A1(new_n2548_), .A2(new_n2549_), .ZN(new_n2630_));
  OAI21_X1  g2438(.A(new_n2551_), .B1(new_n2630_), .B2(new_n2554_), .ZN(new_n2631_));
  XOR2_X1   g2439(.A(new_n2631_), .B(KEYINPUT114), .Z(new_n2632_));
  OR2_X1    g2440(.A1(new_n2629_), .A2(new_n2632_), .ZN(new_n2633_));
  NAND2_X1  g2441(.A1(new_n2629_), .A2(new_n2631_), .ZN(new_n2634_));
  NAND2_X1  g2442(.A1(new_n2633_), .A2(new_n2634_), .ZN(new_n2635_));
  NOR2_X1   g2443(.A1(new_n944_), .A2(new_n918_), .ZN(new_n2636_));
  OR2_X1    g2444(.A1(new_n2635_), .A2(new_n2636_), .ZN(new_n2637_));
  NAND2_X1  g2445(.A1(new_n2635_), .A2(new_n2636_), .ZN(new_n2638_));
  NAND2_X1  g2446(.A1(new_n2637_), .A2(new_n2638_), .ZN(new_n2639_));
  NAND2_X1  g2447(.A1(new_n2571_), .A2(new_n2567_), .ZN(new_n2640_));
  NAND2_X1  g2448(.A1(new_n2639_), .A2(new_n2640_), .ZN(new_n2641_));
  INV_X1    g2449(.A(KEYINPUT115), .ZN(new_n2642_));
  NAND4_X1  g2450(.A1(new_n2637_), .A2(new_n2567_), .A3(new_n2571_), .A4(new_n2638_), .ZN(new_n2643_));
  NAND3_X1  g2451(.A1(new_n2641_), .A2(new_n2642_), .A3(new_n2643_), .ZN(new_n2644_));
  INV_X1    g2452(.A(new_n2643_), .ZN(new_n2645_));
  NAND2_X1  g2453(.A1(new_n2645_), .A2(KEYINPUT115), .ZN(new_n2646_));
  NAND2_X1  g2454(.A1(new_n2644_), .A2(new_n2646_), .ZN(new_n2647_));
  NOR2_X1   g2455(.A1(new_n1093_), .A2(new_n1419_), .ZN(new_n2648_));
  NAND2_X1  g2456(.A1(new_n2647_), .A2(new_n2648_), .ZN(new_n2649_));
  OAI211_X1 g2457(.A(new_n2448_), .B(new_n2577_), .C1(new_n2576_), .C2(new_n2579_), .ZN(new_n2650_));
  NAND2_X1  g2458(.A1(new_n2582_), .A2(new_n2579_), .ZN(new_n2651_));
  AOI21_X1  g2459(.A(new_n2648_), .B1(new_n2641_), .B2(new_n2643_), .ZN(new_n2652_));
  INV_X1    g2460(.A(new_n2652_), .ZN(new_n2653_));
  NAND4_X1  g2461(.A1(new_n2649_), .A2(new_n2650_), .A3(new_n2651_), .A4(new_n2653_), .ZN(new_n2654_));
  INV_X1    g2462(.A(new_n2648_), .ZN(new_n2655_));
  NAND3_X1  g2463(.A1(new_n2644_), .A2(new_n2646_), .A3(new_n2655_), .ZN(new_n2656_));
  NAND3_X1  g2464(.A1(new_n2641_), .A2(new_n2648_), .A3(new_n2643_), .ZN(new_n2657_));
  NAND2_X1  g2465(.A1(new_n2656_), .A2(new_n2657_), .ZN(new_n2658_));
  NAND2_X1  g2466(.A1(new_n2650_), .A2(new_n2651_), .ZN(new_n2659_));
  NAND2_X1  g2467(.A1(new_n2658_), .A2(new_n2659_), .ZN(new_n2660_));
  NAND2_X1  g2468(.A1(new_n2654_), .A2(new_n2660_), .ZN(new_n2661_));
  NOR2_X1   g2469(.A1(new_n799_), .A2(new_n1426_), .ZN(new_n2662_));
  NAND2_X1  g2470(.A1(new_n2661_), .A2(new_n2662_), .ZN(new_n2663_));
  INV_X1    g2471(.A(new_n2662_), .ZN(new_n2664_));
  NAND3_X1  g2472(.A1(new_n2654_), .A2(new_n2660_), .A3(new_n2664_), .ZN(new_n2665_));
  NAND2_X1  g2473(.A1(new_n2663_), .A2(new_n2665_), .ZN(new_n2666_));
  INV_X1    g2474(.A(new_n2587_), .ZN(new_n2667_));
  NAND3_X1  g2475(.A1(new_n2666_), .A2(new_n2667_), .A3(new_n2589_), .ZN(new_n2668_));
  NAND2_X1  g2476(.A1(new_n2589_), .A2(new_n2667_), .ZN(new_n2669_));
  NAND3_X1  g2477(.A1(new_n2669_), .A2(new_n2665_), .A3(new_n2663_), .ZN(new_n2670_));
  NAND2_X1  g2478(.A1(new_n2668_), .A2(new_n2670_), .ZN(new_n2671_));
  NAND3_X1  g2479(.A1(new_n2671_), .A2(G154gat), .A3(G511gat), .ZN(new_n2672_));
  OAI211_X1 g2480(.A(new_n2668_), .B(new_n2670_), .C1(new_n960_), .C2(new_n1438_), .ZN(new_n2673_));
  NAND2_X1  g2481(.A1(new_n2672_), .A2(new_n2673_), .ZN(new_n2674_));
  AOI21_X1  g2482(.A(new_n2591_), .B1(new_n2478_), .B2(new_n2484_), .ZN(new_n2675_));
  NOR2_X1   g2483(.A1(new_n2596_), .A2(new_n2675_), .ZN(new_n2676_));
  NAND2_X1  g2484(.A1(new_n2674_), .A2(new_n2676_), .ZN(new_n2677_));
  INV_X1    g2485(.A(new_n2677_), .ZN(new_n2678_));
  NOR2_X1   g2486(.A1(new_n2674_), .A2(new_n2676_), .ZN(new_n2679_));
  OAI211_X1 g2487(.A(G137gat), .B(G528gat), .C1(new_n2678_), .C2(new_n2679_), .ZN(new_n2680_));
  INV_X1    g2488(.A(new_n2679_), .ZN(new_n2681_));
  NAND2_X1  g2489(.A1(G137gat), .A2(G528gat), .ZN(new_n2682_));
  NAND3_X1  g2490(.A1(new_n2681_), .A2(new_n2682_), .A3(new_n2677_), .ZN(new_n2683_));
  NAND2_X1  g2491(.A1(new_n2680_), .A2(new_n2683_), .ZN(new_n2684_));
  NAND2_X1  g2492(.A1(new_n2606_), .A2(new_n2605_), .ZN(new_n2685_));
  XNOR2_X1  g2493(.A(new_n2684_), .B(new_n2685_), .ZN(new_n2686_));
  XNOR2_X1  g2494(.A(new_n2614_), .B(new_n2686_), .ZN(G6220gat));
  AOI21_X1  g2495(.A(new_n2684_), .B1(new_n2605_), .B2(new_n2606_), .ZN(new_n2688_));
  AOI21_X1  g2496(.A(new_n2688_), .B1(new_n2614_), .B2(new_n2686_), .ZN(new_n2689_));
  NOR2_X1   g2497(.A1(new_n799_), .A2(new_n1438_), .ZN(new_n2690_));
  INV_X1    g2498(.A(new_n2690_), .ZN(new_n2691_));
  NOR2_X1   g2499(.A1(new_n1093_), .A2(new_n1426_), .ZN(new_n2692_));
  INV_X1    g2500(.A(new_n2692_), .ZN(new_n2693_));
  NAND3_X1  g2501(.A1(new_n2640_), .A2(new_n2637_), .A3(new_n2638_), .ZN(new_n2694_));
  OAI21_X1  g2502(.A(new_n2617_), .B1(new_n2619_), .B2(new_n2620_), .ZN(new_n2695_));
  XOR2_X1   g2503(.A(new_n2695_), .B(KEYINPUT117), .Z(new_n2696_));
  NAND2_X1  g2504(.A1(G256gat), .A2(G426gat), .ZN(new_n2697_));
  NAND2_X1  g2505(.A1(new_n2696_), .A2(new_n2697_), .ZN(new_n2698_));
  INV_X1    g2506(.A(new_n2698_), .ZN(new_n2699_));
  NOR2_X1   g2507(.A1(new_n2696_), .A2(new_n2697_), .ZN(new_n2700_));
  NOR2_X1   g2508(.A1(new_n2699_), .A2(new_n2700_), .ZN(new_n2701_));
  NOR2_X1   g2509(.A1(new_n1676_), .A2(new_n768_), .ZN(new_n2702_));
  XOR2_X1   g2510(.A(new_n2701_), .B(new_n2702_), .Z(new_n2703_));
  NOR2_X1   g2511(.A1(new_n2627_), .A2(new_n2628_), .ZN(new_n2704_));
  AOI21_X1  g2512(.A(new_n2621_), .B1(new_n2625_), .B2(new_n2547_), .ZN(new_n2705_));
  NOR2_X1   g2513(.A1(new_n2704_), .A2(new_n2705_), .ZN(new_n2706_));
  OR2_X1    g2514(.A1(new_n2703_), .A2(new_n2706_), .ZN(new_n2707_));
  NOR2_X1   g2515(.A1(new_n1681_), .A2(new_n918_), .ZN(new_n2708_));
  INV_X1    g2516(.A(new_n2708_), .ZN(new_n2709_));
  NAND2_X1  g2517(.A1(new_n2703_), .A2(new_n2706_), .ZN(new_n2710_));
  NAND3_X1  g2518(.A1(new_n2707_), .A2(new_n2709_), .A3(new_n2710_), .ZN(new_n2711_));
  INV_X1    g2519(.A(new_n2711_), .ZN(new_n2712_));
  AOI21_X1  g2520(.A(new_n2709_), .B1(new_n2707_), .B2(new_n2710_), .ZN(new_n2713_));
  NOR2_X1   g2521(.A1(new_n2712_), .A2(new_n2713_), .ZN(new_n2714_));
  NAND2_X1  g2522(.A1(new_n2637_), .A2(new_n2633_), .ZN(new_n2715_));
  NAND2_X1  g2523(.A1(new_n2714_), .A2(new_n2715_), .ZN(new_n2716_));
  NAND2_X1  g2524(.A1(G205gat), .A2(G477gat), .ZN(new_n2717_));
  OAI211_X1 g2525(.A(new_n2637_), .B(new_n2633_), .C1(new_n2712_), .C2(new_n2713_), .ZN(new_n2718_));
  NAND3_X1  g2526(.A1(new_n2716_), .A2(new_n2717_), .A3(new_n2718_), .ZN(new_n2719_));
  INV_X1    g2527(.A(new_n2719_), .ZN(new_n2720_));
  AOI21_X1  g2528(.A(new_n2717_), .B1(new_n2716_), .B2(new_n2718_), .ZN(new_n2721_));
  OAI21_X1  g2529(.A(new_n2694_), .B1(new_n2720_), .B2(new_n2721_), .ZN(new_n2722_));
  NOR2_X1   g2530(.A1(new_n2722_), .A2(new_n2652_), .ZN(new_n2723_));
  INV_X1    g2531(.A(new_n2723_), .ZN(new_n2724_));
  NAND2_X1  g2532(.A1(new_n2656_), .A2(new_n2694_), .ZN(new_n2725_));
  NOR2_X1   g2533(.A1(new_n2720_), .A2(new_n2721_), .ZN(new_n2726_));
  NAND2_X1  g2534(.A1(new_n2725_), .A2(new_n2726_), .ZN(new_n2727_));
  AOI21_X1  g2535(.A(new_n2693_), .B1(new_n2724_), .B2(new_n2727_), .ZN(new_n2728_));
  INV_X1    g2536(.A(new_n2728_), .ZN(new_n2729_));
  INV_X1    g2537(.A(new_n2727_), .ZN(new_n2730_));
  NOR3_X1   g2538(.A1(new_n2730_), .A2(new_n2723_), .A3(new_n2692_), .ZN(new_n2731_));
  INV_X1    g2539(.A(new_n2731_), .ZN(new_n2732_));
  INV_X1    g2540(.A(KEYINPUT118), .ZN(new_n2733_));
  NAND3_X1  g2541(.A1(new_n2729_), .A2(new_n2732_), .A3(new_n2733_), .ZN(new_n2734_));
  OAI21_X1  g2542(.A(KEYINPUT118), .B1(new_n2728_), .B2(new_n2731_), .ZN(new_n2735_));
  OR2_X1    g2543(.A1(new_n2665_), .A2(KEYINPUT116), .ZN(new_n2736_));
  NOR2_X1   g2544(.A1(new_n2658_), .A2(new_n2659_), .ZN(new_n2737_));
  AOI21_X1  g2545(.A(new_n2737_), .B1(new_n2665_), .B2(KEYINPUT116), .ZN(new_n2738_));
  NAND2_X1  g2546(.A1(new_n2736_), .A2(new_n2738_), .ZN(new_n2739_));
  NAND3_X1  g2547(.A1(new_n2734_), .A2(new_n2735_), .A3(new_n2739_), .ZN(new_n2740_));
  NAND2_X1  g2548(.A1(new_n2729_), .A2(new_n2732_), .ZN(new_n2741_));
  NAND4_X1  g2549(.A1(new_n2741_), .A2(KEYINPUT118), .A3(new_n2736_), .A4(new_n2738_), .ZN(new_n2742_));
  AOI21_X1  g2550(.A(new_n2691_), .B1(new_n2740_), .B2(new_n2742_), .ZN(new_n2743_));
  INV_X1    g2551(.A(new_n2743_), .ZN(new_n2744_));
  INV_X1    g2552(.A(KEYINPUT119), .ZN(new_n2745_));
  NAND3_X1  g2553(.A1(new_n2740_), .A2(new_n2742_), .A3(new_n2691_), .ZN(new_n2746_));
  NAND3_X1  g2554(.A1(new_n2744_), .A2(new_n2745_), .A3(new_n2746_), .ZN(new_n2747_));
  INV_X1    g2555(.A(new_n2746_), .ZN(new_n2748_));
  OAI21_X1  g2556(.A(KEYINPUT119), .B1(new_n2748_), .B2(new_n2743_), .ZN(new_n2749_));
  NAND2_X1  g2557(.A1(new_n2673_), .A2(new_n2670_), .ZN(new_n2750_));
  NAND3_X1  g2558(.A1(new_n2747_), .A2(new_n2749_), .A3(new_n2750_), .ZN(new_n2751_));
  AOI21_X1  g2559(.A(new_n2750_), .B1(new_n2744_), .B2(new_n2746_), .ZN(new_n2752_));
  INV_X1    g2560(.A(new_n2752_), .ZN(new_n2753_));
  NAND2_X1  g2561(.A1(new_n2751_), .A2(new_n2753_), .ZN(new_n2754_));
  NOR2_X1   g2562(.A1(new_n960_), .A2(new_n1654_), .ZN(new_n2755_));
  NAND2_X1  g2563(.A1(new_n2754_), .A2(new_n2755_), .ZN(new_n2756_));
  INV_X1    g2564(.A(new_n2755_), .ZN(new_n2757_));
  NAND3_X1  g2565(.A1(new_n2751_), .A2(new_n2757_), .A3(new_n2753_), .ZN(new_n2758_));
  NAND2_X1  g2566(.A1(new_n2756_), .A2(new_n2758_), .ZN(new_n2759_));
  AOI21_X1  g2567(.A(new_n2679_), .B1(new_n2682_), .B2(new_n2677_), .ZN(new_n2760_));
  NAND2_X1  g2568(.A1(new_n2759_), .A2(new_n2760_), .ZN(new_n2761_));
  INV_X1    g2569(.A(new_n2760_), .ZN(new_n2762_));
  NAND3_X1  g2570(.A1(new_n2756_), .A2(new_n2762_), .A3(new_n2758_), .ZN(new_n2763_));
  NAND2_X1  g2571(.A1(new_n2761_), .A2(new_n2763_), .ZN(new_n2764_));
  XNOR2_X1  g2572(.A(new_n2689_), .B(new_n2764_), .ZN(G6230gat));
  NAND3_X1  g2573(.A1(new_n2739_), .A2(new_n2732_), .A3(new_n2729_), .ZN(new_n2766_));
  NAND2_X1  g2574(.A1(new_n2746_), .A2(new_n2766_), .ZN(new_n2767_));
  NOR2_X1   g2575(.A1(new_n1093_), .A2(new_n1438_), .ZN(new_n2768_));
  AND2_X1   g2576(.A1(new_n2711_), .A2(new_n2707_), .ZN(new_n2769_));
  OAI21_X1  g2577(.A(new_n2698_), .B1(new_n2700_), .B2(new_n2702_), .ZN(new_n2770_));
  NAND2_X1  g2578(.A1(G256gat), .A2(G443gat), .ZN(new_n2771_));
  XNOR2_X1  g2579(.A(new_n2770_), .B(new_n2771_), .ZN(new_n2772_));
  NOR2_X1   g2580(.A1(new_n1676_), .A2(new_n918_), .ZN(new_n2773_));
  XNOR2_X1  g2581(.A(new_n2772_), .B(new_n2773_), .ZN(new_n2774_));
  OR2_X1    g2582(.A1(new_n2769_), .A2(new_n2774_), .ZN(new_n2775_));
  NOR2_X1   g2583(.A1(new_n1681_), .A2(new_n1419_), .ZN(new_n2776_));
  INV_X1    g2584(.A(new_n2776_), .ZN(new_n2777_));
  NAND2_X1  g2585(.A1(new_n2769_), .A2(new_n2774_), .ZN(new_n2778_));
  NAND3_X1  g2586(.A1(new_n2775_), .A2(new_n2777_), .A3(new_n2778_), .ZN(new_n2779_));
  INV_X1    g2587(.A(new_n2779_), .ZN(new_n2780_));
  AOI21_X1  g2588(.A(new_n2777_), .B1(new_n2775_), .B2(new_n2778_), .ZN(new_n2781_));
  OAI211_X1 g2589(.A(new_n2716_), .B(new_n2719_), .C1(new_n2780_), .C2(new_n2781_), .ZN(new_n2782_));
  INV_X1    g2590(.A(new_n2781_), .ZN(new_n2783_));
  NAND2_X1  g2591(.A1(new_n2719_), .A2(new_n2716_), .ZN(new_n2784_));
  NAND3_X1  g2592(.A1(new_n2783_), .A2(new_n2784_), .A3(new_n2779_), .ZN(new_n2785_));
  NAND2_X1  g2593(.A1(new_n2782_), .A2(new_n2785_), .ZN(new_n2786_));
  NOR2_X1   g2594(.A1(new_n944_), .A2(new_n1426_), .ZN(new_n2787_));
  XNOR2_X1  g2595(.A(new_n2786_), .B(new_n2787_), .ZN(new_n2788_));
  AOI21_X1  g2596(.A(new_n2730_), .B1(new_n2724_), .B2(new_n2693_), .ZN(new_n2789_));
  NAND2_X1  g2597(.A1(new_n2788_), .A2(new_n2789_), .ZN(new_n2790_));
  INV_X1    g2598(.A(new_n2790_), .ZN(new_n2791_));
  NOR2_X1   g2599(.A1(new_n2788_), .A2(new_n2789_), .ZN(new_n2792_));
  OAI21_X1  g2600(.A(new_n2768_), .B1(new_n2791_), .B2(new_n2792_), .ZN(new_n2793_));
  INV_X1    g2601(.A(new_n2792_), .ZN(new_n2794_));
  INV_X1    g2602(.A(new_n2768_), .ZN(new_n2795_));
  NAND3_X1  g2603(.A1(new_n2794_), .A2(new_n2795_), .A3(new_n2790_), .ZN(new_n2796_));
  AND2_X1   g2604(.A1(new_n2793_), .A2(new_n2796_), .ZN(new_n2797_));
  NAND2_X1  g2605(.A1(new_n2767_), .A2(new_n2797_), .ZN(new_n2798_));
  NAND2_X1  g2606(.A1(new_n2793_), .A2(new_n2796_), .ZN(new_n2799_));
  NAND3_X1  g2607(.A1(new_n2799_), .A2(new_n2746_), .A3(new_n2766_), .ZN(new_n2800_));
  NAND2_X1  g2608(.A1(new_n2798_), .A2(new_n2800_), .ZN(new_n2801_));
  NOR2_X1   g2609(.A1(new_n799_), .A2(new_n1654_), .ZN(new_n2802_));
  NAND2_X1  g2610(.A1(new_n2801_), .A2(new_n2802_), .ZN(new_n2803_));
  OAI211_X1 g2611(.A(new_n2798_), .B(new_n2800_), .C1(new_n799_), .C2(new_n1654_), .ZN(new_n2804_));
  NAND2_X1  g2612(.A1(new_n2803_), .A2(new_n2804_), .ZN(new_n2805_));
  NAND3_X1  g2613(.A1(new_n2805_), .A2(new_n2758_), .A3(new_n2751_), .ZN(new_n2806_));
  OAI21_X1  g2614(.A(new_n2751_), .B1(new_n2752_), .B2(new_n2755_), .ZN(new_n2807_));
  NAND3_X1  g2615(.A1(new_n2807_), .A2(new_n2803_), .A3(new_n2804_), .ZN(new_n2808_));
  AND3_X1   g2616(.A1(new_n2806_), .A2(new_n2808_), .A3(KEYINPUT120), .ZN(new_n2809_));
  AOI21_X1  g2617(.A(KEYINPUT120), .B1(new_n2806_), .B2(new_n2808_), .ZN(new_n2810_));
  NOR2_X1   g2618(.A1(new_n2809_), .A2(new_n2810_), .ZN(new_n2811_));
  OAI21_X1  g2619(.A(new_n2763_), .B1(new_n2689_), .B2(new_n2764_), .ZN(new_n2812_));
  INV_X1    g2620(.A(KEYINPUT121), .ZN(new_n2813_));
  AOI21_X1  g2621(.A(new_n2811_), .B1(new_n2812_), .B2(new_n2813_), .ZN(new_n2814_));
  XNOR2_X1  g2622(.A(new_n2812_), .B(new_n2813_), .ZN(new_n2815_));
  AOI21_X1  g2623(.A(new_n2814_), .B1(new_n2815_), .B2(new_n2811_), .ZN(G6240gat));
  OAI211_X1 g2624(.A(new_n2763_), .B(new_n2808_), .C1(new_n2689_), .C2(new_n2764_), .ZN(new_n2817_));
  NAND2_X1  g2625(.A1(new_n2817_), .A2(new_n2806_), .ZN(new_n2818_));
  NAND2_X1  g2626(.A1(new_n2779_), .A2(new_n2775_), .ZN(new_n2819_));
  NAND2_X1  g2627(.A1(new_n2770_), .A2(new_n2771_), .ZN(new_n2820_));
  OAI21_X1  g2628(.A(new_n2820_), .B1(new_n2772_), .B2(new_n2773_), .ZN(new_n2821_));
  OR3_X1    g2629(.A1(new_n2821_), .A2(new_n1872_), .A3(new_n918_), .ZN(new_n2822_));
  OAI21_X1  g2630(.A(new_n2821_), .B1(new_n1872_), .B2(new_n918_), .ZN(new_n2823_));
  NAND2_X1  g2631(.A1(new_n2822_), .A2(new_n2823_), .ZN(new_n2824_));
  NOR2_X1   g2632(.A1(new_n1676_), .A2(new_n1419_), .ZN(new_n2825_));
  XOR2_X1   g2633(.A(new_n2824_), .B(new_n2825_), .Z(new_n2826_));
  OR2_X1    g2634(.A1(new_n2819_), .A2(new_n2826_), .ZN(new_n2827_));
  NAND2_X1  g2635(.A1(new_n2819_), .A2(new_n2826_), .ZN(new_n2828_));
  NAND2_X1  g2636(.A1(new_n2827_), .A2(new_n2828_), .ZN(new_n2829_));
  NAND3_X1  g2637(.A1(new_n2829_), .A2(G222gat), .A3(G494gat), .ZN(new_n2830_));
  OAI211_X1 g2638(.A(new_n2827_), .B(new_n2828_), .C1(new_n1681_), .C2(new_n1426_), .ZN(new_n2831_));
  AND2_X1   g2639(.A1(new_n2830_), .A2(new_n2831_), .ZN(new_n2832_));
  OAI21_X1  g2640(.A(new_n2785_), .B1(new_n2786_), .B2(new_n2787_), .ZN(new_n2833_));
  XNOR2_X1  g2641(.A(new_n2832_), .B(new_n2833_), .ZN(new_n2834_));
  NOR2_X1   g2642(.A1(new_n944_), .A2(new_n1438_), .ZN(new_n2835_));
  XNOR2_X1  g2643(.A(new_n2834_), .B(new_n2835_), .ZN(new_n2836_));
  AOI21_X1  g2644(.A(new_n2792_), .B1(new_n2795_), .B2(new_n2790_), .ZN(new_n2837_));
  NOR2_X1   g2645(.A1(new_n2836_), .A2(new_n2837_), .ZN(new_n2838_));
  INV_X1    g2646(.A(new_n2838_), .ZN(new_n2839_));
  NOR2_X1   g2647(.A1(new_n1093_), .A2(new_n1654_), .ZN(new_n2840_));
  INV_X1    g2648(.A(new_n2840_), .ZN(new_n2841_));
  NAND2_X1  g2649(.A1(new_n2836_), .A2(new_n2837_), .ZN(new_n2842_));
  AND3_X1   g2650(.A1(new_n2839_), .A2(new_n2841_), .A3(new_n2842_), .ZN(new_n2843_));
  AOI21_X1  g2651(.A(new_n2841_), .B1(new_n2839_), .B2(new_n2842_), .ZN(new_n2844_));
  NOR2_X1   g2652(.A1(new_n2843_), .A2(new_n2844_), .ZN(new_n2845_));
  NAND2_X1  g2653(.A1(new_n2804_), .A2(new_n2798_), .ZN(new_n2846_));
  XNOR2_X1  g2654(.A(new_n2845_), .B(new_n2846_), .ZN(new_n2847_));
  NAND2_X1  g2655(.A1(new_n2818_), .A2(new_n2847_), .ZN(new_n2848_));
  INV_X1    g2656(.A(new_n2847_), .ZN(new_n2849_));
  NAND3_X1  g2657(.A1(new_n2817_), .A2(new_n2806_), .A3(new_n2849_), .ZN(new_n2850_));
  NAND2_X1  g2658(.A1(new_n2848_), .A2(new_n2850_), .ZN(G6250gat));
  AOI21_X1  g2659(.A(new_n2847_), .B1(new_n2811_), .B2(new_n2808_), .ZN(new_n2852_));
  NAND2_X1  g2660(.A1(new_n2817_), .A2(new_n2852_), .ZN(new_n2853_));
  NAND2_X1  g2661(.A1(new_n2853_), .A2(KEYINPUT124), .ZN(new_n2854_));
  NAND2_X1  g2662(.A1(new_n2845_), .A2(new_n2846_), .ZN(new_n2855_));
  INV_X1    g2663(.A(KEYINPUT124), .ZN(new_n2856_));
  NAND3_X1  g2664(.A1(new_n2817_), .A2(new_n2856_), .A3(new_n2852_), .ZN(new_n2857_));
  NAND3_X1  g2665(.A1(new_n2854_), .A2(new_n2855_), .A3(new_n2857_), .ZN(new_n2858_));
  NOR2_X1   g2666(.A1(new_n2843_), .A2(new_n2838_), .ZN(new_n2859_));
  XOR2_X1   g2667(.A(new_n2859_), .B(KEYINPUT123), .Z(new_n2860_));
  NAND2_X1  g2668(.A1(new_n2831_), .A2(new_n2828_), .ZN(new_n2861_));
  OAI21_X1  g2669(.A(new_n2823_), .B1(new_n2824_), .B2(new_n2825_), .ZN(new_n2862_));
  OR3_X1    g2670(.A1(new_n2862_), .A2(new_n1872_), .A3(new_n1419_), .ZN(new_n2863_));
  OAI21_X1  g2671(.A(new_n2862_), .B1(new_n1872_), .B2(new_n1419_), .ZN(new_n2864_));
  NAND2_X1  g2672(.A1(new_n2863_), .A2(new_n2864_), .ZN(new_n2865_));
  NOR2_X1   g2673(.A1(new_n1676_), .A2(new_n1426_), .ZN(new_n2866_));
  XOR2_X1   g2674(.A(new_n2865_), .B(new_n2866_), .Z(new_n2867_));
  XNOR2_X1  g2675(.A(new_n2861_), .B(new_n2867_), .ZN(new_n2868_));
  XOR2_X1   g2676(.A(new_n2868_), .B(KEYINPUT122), .Z(new_n2869_));
  NOR2_X1   g2677(.A1(new_n1681_), .A2(new_n1438_), .ZN(new_n2870_));
  OR2_X1    g2678(.A1(new_n2869_), .A2(new_n2870_), .ZN(new_n2871_));
  NAND2_X1  g2679(.A1(new_n2869_), .A2(new_n2870_), .ZN(new_n2872_));
  NAND2_X1  g2680(.A1(new_n2871_), .A2(new_n2872_), .ZN(new_n2873_));
  NAND2_X1  g2681(.A1(new_n2832_), .A2(new_n2833_), .ZN(new_n2874_));
  OAI21_X1  g2682(.A(new_n2874_), .B1(new_n2834_), .B2(new_n2835_), .ZN(new_n2875_));
  XNOR2_X1  g2683(.A(new_n2873_), .B(new_n2875_), .ZN(new_n2876_));
  NAND2_X1  g2684(.A1(G205gat), .A2(G528gat), .ZN(new_n2877_));
  XNOR2_X1  g2685(.A(new_n2876_), .B(new_n2877_), .ZN(new_n2878_));
  OR2_X1    g2686(.A1(new_n2860_), .A2(new_n2878_), .ZN(new_n2879_));
  NAND2_X1  g2687(.A1(new_n2860_), .A2(new_n2878_), .ZN(new_n2880_));
  AND2_X1   g2688(.A1(new_n2879_), .A2(new_n2880_), .ZN(new_n2881_));
  NAND2_X1  g2689(.A1(new_n2858_), .A2(new_n2881_), .ZN(new_n2882_));
  NAND2_X1  g2690(.A1(new_n2850_), .A2(new_n2855_), .ZN(new_n2883_));
  OAI21_X1  g2691(.A(new_n2882_), .B1(new_n2881_), .B2(new_n2883_), .ZN(G6260gat));
  NAND3_X1  g2692(.A1(new_n2850_), .A2(new_n2855_), .A3(new_n2879_), .ZN(new_n2885_));
  NAND2_X1  g2693(.A1(new_n2885_), .A2(new_n2880_), .ZN(new_n2886_));
  NAND2_X1  g2694(.A1(new_n2861_), .A2(new_n2867_), .ZN(new_n2887_));
  NAND2_X1  g2695(.A1(new_n2871_), .A2(new_n2887_), .ZN(new_n2888_));
  OAI21_X1  g2696(.A(new_n2864_), .B1(new_n2865_), .B2(new_n2866_), .ZN(new_n2889_));
  OR3_X1    g2697(.A1(new_n2889_), .A2(new_n1872_), .A3(new_n1426_), .ZN(new_n2890_));
  OAI21_X1  g2698(.A(new_n2889_), .B1(new_n1872_), .B2(new_n1426_), .ZN(new_n2891_));
  NAND2_X1  g2699(.A1(new_n2890_), .A2(new_n2891_), .ZN(new_n2892_));
  XOR2_X1   g2700(.A(new_n2892_), .B(KEYINPUT125), .Z(new_n2893_));
  NAND2_X1  g2701(.A1(G239gat), .A2(G511gat), .ZN(new_n2894_));
  NAND2_X1  g2702(.A1(new_n2893_), .A2(new_n2894_), .ZN(new_n2895_));
  INV_X1    g2703(.A(new_n2895_), .ZN(new_n2896_));
  NOR2_X1   g2704(.A1(new_n2893_), .A2(new_n2894_), .ZN(new_n2897_));
  NOR2_X1   g2705(.A1(new_n2896_), .A2(new_n2897_), .ZN(new_n2898_));
  NAND2_X1  g2706(.A1(new_n2888_), .A2(new_n2898_), .ZN(new_n2899_));
  INV_X1    g2707(.A(new_n2899_), .ZN(new_n2900_));
  NOR2_X1   g2708(.A1(new_n1681_), .A2(new_n1654_), .ZN(new_n2901_));
  NOR2_X1   g2709(.A1(new_n2888_), .A2(new_n2898_), .ZN(new_n2902_));
  OR3_X1    g2710(.A1(new_n2900_), .A2(new_n2901_), .A3(new_n2902_), .ZN(new_n2903_));
  OAI21_X1  g2711(.A(new_n2901_), .B1(new_n2900_), .B2(new_n2902_), .ZN(new_n2904_));
  AND2_X1   g2712(.A1(new_n2903_), .A2(new_n2904_), .ZN(new_n2905_));
  NAND2_X1  g2713(.A1(new_n2876_), .A2(new_n2877_), .ZN(new_n2906_));
  NAND3_X1  g2714(.A1(new_n2871_), .A2(new_n2875_), .A3(new_n2872_), .ZN(new_n2907_));
  NAND2_X1  g2715(.A1(new_n2906_), .A2(new_n2907_), .ZN(new_n2908_));
  NOR2_X1   g2716(.A1(new_n2905_), .A2(new_n2908_), .ZN(new_n2909_));
  INV_X1    g2717(.A(new_n2909_), .ZN(new_n2910_));
  NAND2_X1  g2718(.A1(new_n2905_), .A2(new_n2908_), .ZN(new_n2911_));
  AND2_X1   g2719(.A1(new_n2910_), .A2(new_n2911_), .ZN(new_n2912_));
  XOR2_X1   g2720(.A(new_n2886_), .B(new_n2912_), .Z(G6270gat));
  NAND2_X1  g2721(.A1(new_n2903_), .A2(new_n2899_), .ZN(new_n2914_));
  INV_X1    g2722(.A(new_n2914_), .ZN(new_n2915_));
  NOR2_X1   g2723(.A1(new_n2896_), .A2(KEYINPUT126), .ZN(new_n2916_));
  INV_X1    g2724(.A(KEYINPUT126), .ZN(new_n2917_));
  OAI21_X1  g2725(.A(new_n2891_), .B1(new_n2895_), .B2(new_n2917_), .ZN(new_n2918_));
  NOR2_X1   g2726(.A1(new_n2916_), .A2(new_n2918_), .ZN(new_n2919_));
  NOR2_X1   g2727(.A1(new_n1872_), .A2(new_n1438_), .ZN(new_n2920_));
  AND2_X1   g2728(.A1(new_n2919_), .A2(new_n2920_), .ZN(new_n2921_));
  NOR2_X1   g2729(.A1(new_n2919_), .A2(new_n2920_), .ZN(new_n2922_));
  NOR2_X1   g2730(.A1(new_n2921_), .A2(new_n2922_), .ZN(new_n2923_));
  NOR2_X1   g2731(.A1(new_n1676_), .A2(new_n1654_), .ZN(new_n2924_));
  XNOR2_X1  g2732(.A(new_n2923_), .B(new_n2924_), .ZN(new_n2925_));
  INV_X1    g2733(.A(new_n2925_), .ZN(new_n2926_));
  NOR2_X1   g2734(.A1(new_n2915_), .A2(new_n2926_), .ZN(new_n2927_));
  INV_X1    g2735(.A(new_n2927_), .ZN(new_n2928_));
  NAND2_X1  g2736(.A1(new_n2915_), .A2(new_n2926_), .ZN(new_n2929_));
  AND2_X1   g2737(.A1(new_n2928_), .A2(new_n2929_), .ZN(new_n2930_));
  NAND3_X1  g2738(.A1(new_n2885_), .A2(new_n2880_), .A3(new_n2912_), .ZN(new_n2931_));
  NAND2_X1  g2739(.A1(new_n2931_), .A2(new_n2911_), .ZN(new_n2932_));
  NAND2_X1  g2740(.A1(new_n2879_), .A2(new_n2911_), .ZN(new_n2933_));
  AOI21_X1  g2741(.A(new_n2933_), .B1(new_n2858_), .B2(new_n2881_), .ZN(new_n2934_));
  NAND2_X1  g2742(.A1(new_n2930_), .A2(new_n2910_), .ZN(new_n2935_));
  OAI22_X1  g2743(.A1(new_n2930_), .A2(new_n2932_), .B1(new_n2934_), .B2(new_n2935_), .ZN(G6280gat));
  OAI21_X1  g2744(.A(new_n2928_), .B1(new_n2934_), .B2(new_n2935_), .ZN(new_n2937_));
  INV_X1    g2745(.A(new_n2922_), .ZN(new_n2938_));
  OAI21_X1  g2746(.A(new_n2938_), .B1(new_n2921_), .B2(new_n2924_), .ZN(new_n2939_));
  OR2_X1    g2747(.A1(new_n2939_), .A2(KEYINPUT127), .ZN(new_n2940_));
  NOR2_X1   g2748(.A1(new_n1872_), .A2(new_n1654_), .ZN(new_n2941_));
  NAND2_X1  g2749(.A1(new_n2939_), .A2(KEYINPUT127), .ZN(new_n2942_));
  AND3_X1   g2750(.A1(new_n2940_), .A2(new_n2941_), .A3(new_n2942_), .ZN(new_n2943_));
  AOI21_X1  g2751(.A(new_n2941_), .B1(new_n2940_), .B2(new_n2942_), .ZN(new_n2944_));
  NOR2_X1   g2752(.A1(new_n2943_), .A2(new_n2944_), .ZN(new_n2945_));
  INV_X1    g2753(.A(new_n2945_), .ZN(new_n2946_));
  INV_X1    g2754(.A(new_n2941_), .ZN(new_n2947_));
  AOI22_X1  g2755(.A1(new_n2937_), .A2(new_n2946_), .B1(new_n2947_), .B2(new_n2939_), .ZN(G6287gat));
  NAND2_X1  g2756(.A1(new_n2932_), .A2(new_n2929_), .ZN(new_n2949_));
  NOR2_X1   g2757(.A1(new_n2945_), .A2(new_n2927_), .ZN(new_n2950_));
  AOI22_X1  g2758(.A1(new_n2937_), .A2(new_n2945_), .B1(new_n2949_), .B2(new_n2950_), .ZN(G6288gat));
endmodule


