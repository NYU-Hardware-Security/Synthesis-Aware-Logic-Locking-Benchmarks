//Secret key is'0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_c2670" written by ABC on Wed Nov 16 09:33:23 2022

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14,
    G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32,
    G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52,
    G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68,
    G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101,
    G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115,
    G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129,
    G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169,
    G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189,
    G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
    G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213,
    G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248,
    G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264,
    G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276,
    G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860, G868,
    G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981,
    G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096,
    G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446,
    G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445_, new_n447_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n457_, new_n458_, new_n459_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n528_, new_n529_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n541_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n581_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_;
  XOR2_X1   g000(.A(KEYINPUT0), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT1), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  INV_X1    g010(.A(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT3), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT4), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445_));
  XOR2_X1   g020(.A(new_n445_), .B(KEYINPUT5), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447_));
  XNOR2_X1  g022(.A(new_n447_), .B(KEYINPUT6), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n451_));
  XNOR2_X1  g026(.A(new_n451_), .B(KEYINPUT7), .ZN(new_n452_));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453_));
  INV_X1    g028(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g029(.A1(new_n452_), .A2(new_n454_), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452_), .A2(G567), .ZN(new_n457_));
  INV_X1    g032(.A(G2106), .ZN(new_n458_));
  OAI21_X1  g033(.A(new_n457_), .B1(new_n458_), .B2(new_n453_), .ZN(new_n459_));
  INV_X1    g034(.A(new_n459_), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT10), .ZN(new_n461_));
  AND2_X1   g036(.A1(KEYINPUT9), .A2(G2104), .ZN(new_n462_));
  NOR2_X1   g037(.A1(KEYINPUT9), .A2(G2104), .ZN(new_n463_));
  NOR2_X1   g038(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND2_X1   g039(.A1(G125), .A2(G2105), .ZN(new_n465_));
  AOI21_X1  g040(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OR2_X1    g041(.A1(KEYINPUT9), .A2(G2104), .ZN(new_n467_));
  NAND2_X1  g042(.A1(KEYINPUT9), .A2(G2104), .ZN(new_n468_));
  AND4_X1   g043(.A1(new_n461_), .A2(new_n467_), .A3(new_n468_), .A4(new_n465_), .ZN(new_n469_));
  NOR2_X1   g044(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g045(.A(G2105), .ZN(new_n471_));
  NAND2_X1  g046(.A1(new_n471_), .A2(KEYINPUT8), .ZN(new_n472_));
  INV_X1    g047(.A(KEYINPUT8), .ZN(new_n473_));
  NAND2_X1  g048(.A1(new_n473_), .A2(G2105), .ZN(new_n474_));
  NAND4_X1  g049(.A1(new_n472_), .A2(new_n474_), .A3(G101), .A4(G2104), .ZN(new_n475_));
  NAND3_X1  g050(.A1(G113), .A2(G2104), .A3(G2105), .ZN(new_n476_));
  NAND4_X1  g051(.A1(new_n467_), .A2(new_n472_), .A3(new_n474_), .A4(new_n468_), .ZN(new_n477_));
  INV_X1    g052(.A(G137), .ZN(new_n478_));
  OAI211_X1 g053(.A(new_n475_), .B(new_n476_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g054(.A1(new_n470_), .A2(new_n479_), .ZN(G160));
  XNOR2_X1  g055(.A(KEYINPUT8), .B(G2105), .ZN(new_n481_));
  AND2_X1   g056(.A1(new_n481_), .A2(G2104), .ZN(new_n482_));
  AND4_X1   g057(.A1(new_n467_), .A2(new_n472_), .A3(new_n474_), .A4(new_n468_), .ZN(new_n483_));
  AOI22_X1  g058(.A1(new_n482_), .A2(G100), .B1(new_n483_), .B2(G136), .ZN(new_n484_));
  AOI22_X1  g059(.A1(new_n464_), .A2(G124), .B1(G112), .B2(G2104), .ZN(new_n485_));
  OAI21_X1  g060(.A(new_n484_), .B1(new_n471_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g061(.A(new_n486_), .B(KEYINPUT11), .ZN(new_n487_));
  XNOR2_X1  g062(.A(new_n487_), .B(KEYINPUT12), .ZN(G162));
  AND3_X1   g063(.A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n489_));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490_));
  AOI21_X1  g065(.A(new_n489_), .B1(new_n464_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g066(.A1(new_n464_), .A2(new_n481_), .A3(G138), .ZN(new_n492_));
  NAND3_X1  g067(.A1(new_n481_), .A2(G102), .A3(G2104), .ZN(new_n493_));
  NAND3_X1  g068(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  XOR2_X1   g069(.A(new_n494_), .B(KEYINPUT13), .Z(G164));
  INV_X1    g070(.A(G651), .ZN(new_n496_));
  NAND3_X1  g071(.A1(new_n496_), .A2(G50), .A3(G543), .ZN(new_n497_));
  INV_X1    g072(.A(KEYINPUT14), .ZN(new_n498_));
  XNOR2_X1  g073(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  NOR2_X1   g074(.A1(G543), .A2(G651), .ZN(new_n500_));
  NAND2_X1  g075(.A1(new_n500_), .A2(G88), .ZN(new_n501_));
  INV_X1    g076(.A(G543), .ZN(new_n502_));
  NOR2_X1   g077(.A1(new_n502_), .A2(G75), .ZN(new_n503_));
  OAI21_X1  g078(.A(G651), .B1(G62), .B2(G543), .ZN(new_n504_));
  OAI211_X1 g079(.A(new_n499_), .B(new_n501_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g080(.A(new_n505_), .B(KEYINPUT15), .ZN(G166));
  NAND3_X1  g081(.A1(new_n496_), .A2(G51), .A3(G543), .ZN(new_n507_));
  XOR2_X1   g082(.A(new_n507_), .B(KEYINPUT17), .Z(new_n508_));
  NOR2_X1   g083(.A1(new_n502_), .A2(G76), .ZN(new_n509_));
  OAI21_X1  g084(.A(G651), .B1(G63), .B2(G543), .ZN(new_n510_));
  OAI21_X1  g085(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g086(.A1(new_n500_), .A2(G89), .ZN(new_n512_));
  XOR2_X1   g087(.A(new_n512_), .B(KEYINPUT16), .Z(new_n513_));
  NOR2_X1   g088(.A1(new_n511_), .A2(new_n513_), .ZN(G168));
  AOI21_X1  g089(.A(new_n496_), .B1(G64), .B2(new_n502_), .ZN(new_n515_));
  INV_X1    g090(.A(G77), .ZN(new_n516_));
  OAI21_X1  g091(.A(new_n515_), .B1(new_n516_), .B2(new_n502_), .ZN(new_n517_));
  AOI21_X1  g092(.A(G651), .B1(new_n502_), .B2(G90), .ZN(new_n518_));
  INV_X1    g093(.A(G52), .ZN(new_n519_));
  OAI21_X1  g094(.A(new_n518_), .B1(new_n519_), .B2(new_n502_), .ZN(new_n520_));
  NAND2_X1  g095(.A1(new_n517_), .A2(new_n520_), .ZN(G171));
  OR2_X1    g096(.A1(G56), .A2(G543), .ZN(new_n522_));
  OAI211_X1 g097(.A(new_n522_), .B(G651), .C1(G68), .C2(new_n502_), .ZN(new_n523_));
  OR2_X1    g098(.A1(G81), .A2(G543), .ZN(new_n524_));
  OAI211_X1 g099(.A(new_n524_), .B(new_n496_), .C1(G43), .C2(new_n502_), .ZN(new_n525_));
  NAND3_X1  g100(.A1(new_n523_), .A2(new_n525_), .A3(G860), .ZN(G153));
  NAND4_X1  g101(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g102(.A1(G1), .A2(G3), .ZN(new_n528_));
  NAND4_X1  g103(.A1(G319), .A2(G483), .A3(G661), .A4(new_n528_), .ZN(new_n529_));
  XOR2_X1   g104(.A(new_n529_), .B(KEYINPUT18), .Z(G188));
  AOI21_X1  g105(.A(new_n496_), .B1(G65), .B2(new_n502_), .ZN(new_n531_));
  INV_X1    g106(.A(G78), .ZN(new_n532_));
  OAI21_X1  g107(.A(new_n531_), .B1(new_n532_), .B2(new_n502_), .ZN(new_n533_));
  AOI21_X1  g108(.A(G651), .B1(new_n502_), .B2(G91), .ZN(new_n534_));
  INV_X1    g109(.A(G53), .ZN(new_n535_));
  OAI21_X1  g110(.A(new_n534_), .B1(new_n535_), .B2(new_n502_), .ZN(new_n536_));
  NAND2_X1  g111(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g112(.A(new_n537_), .ZN(G299));
  INV_X1    g113(.A(G171), .ZN(G301));
  INV_X1    g114(.A(G168), .ZN(G286));
  INV_X1    g115(.A(KEYINPUT15), .ZN(new_n541_));
  XNOR2_X1  g116(.A(new_n505_), .B(new_n541_), .ZN(G303));
  NAND2_X1  g117(.A1(G49), .A2(G543), .ZN(new_n543_));
  INV_X1    g118(.A(G87), .ZN(new_n544_));
  OAI211_X1 g119(.A(new_n543_), .B(new_n496_), .C1(new_n544_), .C2(G543), .ZN(new_n545_));
  INV_X1    g120(.A(G74), .ZN(new_n546_));
  NAND3_X1  g121(.A1(new_n546_), .A2(G543), .A3(G651), .ZN(new_n547_));
  NAND2_X1  g122(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g123(.A(KEYINPUT19), .ZN(new_n549_));
  XNOR2_X1  g124(.A(new_n548_), .B(new_n549_), .ZN(G288));
  AOI21_X1  g125(.A(new_n496_), .B1(G61), .B2(new_n502_), .ZN(new_n551_));
  INV_X1    g126(.A(G73), .ZN(new_n552_));
  OAI21_X1  g127(.A(new_n551_), .B1(new_n552_), .B2(new_n502_), .ZN(new_n553_));
  AOI21_X1  g128(.A(G651), .B1(new_n502_), .B2(G86), .ZN(new_n554_));
  INV_X1    g129(.A(G48), .ZN(new_n555_));
  OAI21_X1  g130(.A(new_n554_), .B1(new_n555_), .B2(new_n502_), .ZN(new_n556_));
  NAND2_X1  g131(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g132(.A(new_n557_), .ZN(G305));
  NAND3_X1  g133(.A1(new_n496_), .A2(G47), .A3(G543), .ZN(new_n559_));
  XOR2_X1   g134(.A(new_n559_), .B(KEYINPUT21), .Z(new_n560_));
  NAND2_X1  g135(.A1(new_n500_), .A2(G85), .ZN(new_n561_));
  XNOR2_X1  g136(.A(new_n561_), .B(KEYINPUT20), .ZN(new_n562_));
  NAND3_X1  g137(.A1(G72), .A2(G543), .A3(G651), .ZN(new_n563_));
  NAND3_X1  g138(.A1(new_n502_), .A2(G60), .A3(G651), .ZN(new_n564_));
  XNOR2_X1  g139(.A(new_n564_), .B(KEYINPUT22), .ZN(new_n565_));
  NAND4_X1  g140(.A1(new_n560_), .A2(new_n562_), .A3(new_n563_), .A4(new_n565_), .ZN(G290));
  NAND2_X1  g141(.A1(new_n500_), .A2(G92), .ZN(new_n567_));
  NOR2_X1   g142(.A1(new_n502_), .A2(G79), .ZN(new_n568_));
  OAI21_X1  g143(.A(G651), .B1(G66), .B2(G543), .ZN(new_n569_));
  OAI21_X1  g144(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n571_));
  NAND2_X1  g146(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g147(.A(new_n567_), .B(KEYINPUT23), .C1(new_n568_), .C2(new_n569_), .ZN(new_n573_));
  NAND2_X1  g148(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g149(.A1(new_n496_), .A2(G54), .A3(G543), .ZN(new_n575_));
  NAND2_X1  g150(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g151(.A(new_n576_), .B(KEYINPUT24), .ZN(new_n577_));
  INV_X1    g152(.A(new_n577_), .ZN(new_n578_));
  MUX2_X1   g153(.A(new_n578_), .B(G301), .S(G868), .Z(G284));
  XNOR2_X1  g154(.A(G284), .B(KEYINPUT25), .ZN(G321));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G868), .ZN(new_n581_));
  MUX2_X1   g156(.A(G286), .B(G299), .S(new_n581_), .Z(G297));
  MUX2_X1   g157(.A(G286), .B(G299), .S(new_n581_), .Z(G280));
  INV_X1    g158(.A(G559), .ZN(new_n584_));
  AOI21_X1  g159(.A(G860), .B1(new_n584_), .B2(KEYINPUT27), .ZN(new_n585_));
  OAI21_X1  g160(.A(new_n585_), .B1(KEYINPUT27), .B2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g161(.A1(new_n577_), .A2(new_n586_), .ZN(G148));
  INV_X1    g162(.A(new_n576_), .ZN(new_n588_));
  NAND2_X1  g163(.A1(new_n588_), .A2(new_n584_), .ZN(new_n589_));
  NAND2_X1  g164(.A1(new_n523_), .A2(new_n525_), .ZN(new_n590_));
  MUX2_X1   g165(.A(new_n589_), .B(new_n590_), .S(new_n581_), .Z(G282));
  MUX2_X1   g166(.A(new_n589_), .B(new_n590_), .S(new_n581_), .Z(G323));
  NAND2_X1  g167(.A1(new_n482_), .A2(G99), .ZN(new_n593_));
  NAND2_X1  g168(.A1(new_n467_), .A2(new_n468_), .ZN(new_n594_));
  NOR2_X1   g169(.A1(new_n594_), .A2(new_n471_), .ZN(new_n595_));
  NAND2_X1  g170(.A1(new_n595_), .A2(G123), .ZN(new_n596_));
  NAND2_X1  g171(.A1(new_n483_), .A2(G135), .ZN(new_n597_));
  NAND3_X1  g172(.A1(G111), .A2(G2104), .A3(G2105), .ZN(new_n598_));
  XOR2_X1   g173(.A(new_n598_), .B(KEYINPUT28), .Z(new_n599_));
  NAND4_X1  g174(.A1(new_n593_), .A2(new_n596_), .A3(new_n597_), .A4(new_n599_), .ZN(new_n600_));
  XOR2_X1   g175(.A(new_n600_), .B(KEYINPUT29), .Z(new_n601_));
  OR2_X1    g176(.A1(new_n601_), .A2(G2096), .ZN(new_n602_));
  NAND2_X1  g177(.A1(new_n601_), .A2(G2096), .ZN(new_n603_));
  INV_X1    g178(.A(KEYINPUT9), .ZN(new_n604_));
  OAI21_X1  g179(.A(new_n482_), .B1(KEYINPUT8), .B2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g180(.A(new_n605_), .B(G2100), .Z(new_n606_));
  NAND3_X1  g181(.A1(new_n602_), .A2(new_n603_), .A3(new_n606_), .ZN(G156));
  XNOR2_X1  g182(.A(G1341), .B(G1348), .ZN(new_n608_));
  XNOR2_X1  g183(.A(KEYINPUT33), .B(G2454), .ZN(new_n609_));
  XNOR2_X1  g184(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g185(.A(new_n610_), .ZN(new_n611_));
  XOR2_X1   g186(.A(G2427), .B(G2430), .Z(new_n612_));
  XOR2_X1   g187(.A(G2435), .B(G2438), .Z(new_n613_));
  OR2_X1    g188(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g189(.A(G2443), .B(G2446), .ZN(new_n615_));
  NOR2_X1   g190(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g191(.A(new_n616_), .B(KEYINPUT31), .ZN(new_n617_));
  NAND2_X1  g192(.A1(new_n612_), .A2(new_n613_), .ZN(new_n618_));
  NOR2_X1   g193(.A1(new_n618_), .A2(new_n615_), .ZN(new_n619_));
  XNOR2_X1  g194(.A(new_n619_), .B(KEYINPUT30), .ZN(new_n620_));
  NAND3_X1  g195(.A1(new_n614_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n621_));
  NAND3_X1  g196(.A1(new_n617_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g197(.A1(new_n622_), .A2(KEYINPUT32), .ZN(new_n623_));
  INV_X1    g198(.A(G2451), .ZN(new_n624_));
  INV_X1    g199(.A(KEYINPUT32), .ZN(new_n625_));
  NAND4_X1  g200(.A1(new_n617_), .A2(new_n625_), .A3(new_n620_), .A4(new_n621_), .ZN(new_n626_));
  NAND3_X1  g201(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g202(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g203(.A(new_n624_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n629_));
  OAI21_X1  g204(.A(new_n611_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g205(.A(new_n629_), .ZN(new_n631_));
  NAND3_X1  g206(.A1(new_n631_), .A2(new_n627_), .A3(new_n610_), .ZN(new_n632_));
  NAND3_X1  g207(.A1(new_n630_), .A2(new_n632_), .A3(G14), .ZN(new_n633_));
  INV_X1    g208(.A(new_n633_), .ZN(G401));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635_));
  XOR2_X1   g210(.A(G2072), .B(G2078), .Z(new_n636_));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637_));
  OR2_X1    g212(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g213(.A(KEYINPUT34), .ZN(new_n639_));
  NAND2_X1  g214(.A1(new_n636_), .A2(new_n637_), .ZN(new_n640_));
  NAND3_X1  g215(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g216(.A1(new_n641_), .A2(KEYINPUT35), .ZN(new_n642_));
  INV_X1    g217(.A(KEYINPUT35), .ZN(new_n643_));
  NAND2_X1  g218(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g219(.A(new_n635_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g220(.A(new_n645_), .B1(new_n635_), .B2(new_n642_), .ZN(new_n646_));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647_));
  XOR2_X1   g222(.A(new_n646_), .B(new_n647_), .Z(new_n648_));
  XNOR2_X1  g223(.A(KEYINPUT36), .B(KEYINPUT37), .ZN(new_n649_));
  XNOR2_X1  g224(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g225(.A(new_n650_), .ZN(G227));
  XNOR2_X1  g226(.A(G1981), .B(G1986), .ZN(new_n652_));
  XNOR2_X1  g227(.A(new_n652_), .B(KEYINPUT42), .ZN(new_n653_));
  XNOR2_X1  g228(.A(G1961), .B(G1966), .ZN(new_n654_));
  INV_X1    g229(.A(KEYINPUT38), .ZN(new_n655_));
  XNOR2_X1  g230(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657_));
  NAND2_X1  g232(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659_));
  XNOR2_X1  g234(.A(new_n659_), .B(KEYINPUT39), .ZN(new_n660_));
  NOR2_X1   g235(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g236(.A(KEYINPUT40), .ZN(new_n662_));
  XNOR2_X1  g237(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  INV_X1    g238(.A(KEYINPUT41), .ZN(new_n664_));
  NAND2_X1  g239(.A1(new_n658_), .A2(new_n660_), .ZN(new_n665_));
  NOR2_X1   g240(.A1(new_n656_), .A2(new_n657_), .ZN(new_n666_));
  MUX2_X1   g241(.A(new_n665_), .B(new_n660_), .S(new_n666_), .Z(new_n667_));
  NAND3_X1  g242(.A1(new_n663_), .A2(new_n664_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g243(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g244(.A(new_n664_), .B1(new_n663_), .B2(new_n667_), .ZN(new_n670_));
  OAI21_X1  g245(.A(new_n653_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g246(.A(new_n670_), .ZN(new_n672_));
  INV_X1    g247(.A(new_n653_), .ZN(new_n673_));
  NAND3_X1  g248(.A1(new_n672_), .A2(new_n673_), .A3(new_n668_), .ZN(new_n674_));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675_));
  AND3_X1   g250(.A1(new_n671_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g251(.A(new_n675_), .B1(new_n671_), .B2(new_n674_), .ZN(new_n677_));
  NOR2_X1   g252(.A1(new_n676_), .A2(new_n677_), .ZN(G229));
  NAND2_X1  g253(.A1(G166), .A2(G16), .ZN(new_n679_));
  OAI21_X1  g254(.A(new_n679_), .B1(G16), .B2(G22), .ZN(new_n680_));
  XNOR2_X1  g255(.A(KEYINPUT71), .B(G1971), .ZN(new_n681_));
  AND2_X1   g256(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g257(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  INV_X1    g258(.A(G29), .ZN(new_n684_));
  AND2_X1   g259(.A1(KEYINPUT58), .A2(G32), .ZN(new_n685_));
  NOR2_X1   g260(.A1(KEYINPUT58), .A2(G32), .ZN(new_n686_));
  OAI21_X1  g261(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g262(.A(new_n687_), .B(KEYINPUT59), .ZN(new_n688_));
  NAND2_X1  g263(.A1(new_n483_), .A2(G141), .ZN(new_n689_));
  XNOR2_X1  g264(.A(new_n689_), .B(KEYINPUT60), .ZN(new_n690_));
  NAND2_X1  g265(.A1(G117), .A2(G2104), .ZN(new_n691_));
  INV_X1    g266(.A(G129), .ZN(new_n692_));
  OAI21_X1  g267(.A(new_n691_), .B1(new_n594_), .B2(new_n692_), .ZN(new_n693_));
  AOI22_X1  g268(.A1(G2105), .A2(new_n693_), .B1(new_n482_), .B2(G105), .ZN(new_n694_));
  NAND2_X1  g269(.A1(new_n690_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g270(.A(new_n688_), .B1(new_n695_), .B2(G29), .ZN(new_n696_));
  XOR2_X1   g271(.A(KEYINPUT61), .B(G1996), .Z(new_n697_));
  NOR2_X1   g272(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g273(.A1(new_n682_), .A2(new_n683_), .A3(new_n698_), .ZN(new_n699_));
  AOI22_X1  g274(.A1(new_n464_), .A2(G119), .B1(G107), .B2(G2104), .ZN(new_n700_));
  NOR2_X1   g275(.A1(new_n700_), .A2(new_n471_), .ZN(new_n701_));
  NAND2_X1  g276(.A1(new_n481_), .A2(G2104), .ZN(new_n702_));
  INV_X1    g277(.A(G95), .ZN(new_n703_));
  INV_X1    g278(.A(G131), .ZN(new_n704_));
  OAI22_X1  g279(.A1(new_n702_), .A2(new_n703_), .B1(new_n477_), .B2(new_n704_), .ZN(new_n705_));
  OR3_X1    g280(.A1(new_n701_), .A2(new_n705_), .A3(KEYINPUT73), .ZN(new_n706_));
  OAI21_X1  g281(.A(KEYINPUT73), .B1(new_n701_), .B2(new_n705_), .ZN(new_n707_));
  NAND2_X1  g282(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  MUX2_X1   g283(.A(G25), .B(new_n708_), .S(G29), .Z(new_n709_));
  NOR2_X1   g284(.A1(new_n709_), .A2(G1991), .ZN(new_n710_));
  OR2_X1    g285(.A1(KEYINPUT72), .A2(G23), .ZN(new_n711_));
  NAND2_X1  g286(.A1(KEYINPUT72), .A2(G23), .ZN(new_n712_));
  AOI21_X1  g287(.A(G16), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g288(.A(new_n713_), .B1(G288), .B2(G16), .ZN(new_n714_));
  XOR2_X1   g289(.A(new_n714_), .B(G1976), .Z(new_n715_));
  INV_X1    g290(.A(G16), .ZN(new_n716_));
  AND2_X1   g291(.A1(new_n716_), .A2(G24), .ZN(new_n717_));
  AOI21_X1  g292(.A(new_n717_), .B1(G290), .B2(G16), .ZN(new_n718_));
  INV_X1    g293(.A(G1986), .ZN(new_n719_));
  OAI22_X1  g294(.A1(new_n601_), .A2(new_n684_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g295(.A1(new_n710_), .A2(new_n715_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g296(.A1(new_n482_), .A2(G103), .ZN(new_n722_));
  NAND2_X1  g297(.A1(new_n595_), .A2(G127), .ZN(new_n723_));
  NAND2_X1  g298(.A1(new_n483_), .A2(G139), .ZN(new_n724_));
  NAND3_X1  g299(.A1(G115), .A2(G2104), .A3(G2105), .ZN(new_n725_));
  XNOR2_X1  g300(.A(new_n725_), .B(KEYINPUT56), .ZN(new_n726_));
  NAND4_X1  g301(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .A4(new_n726_), .ZN(new_n727_));
  MUX2_X1   g302(.A(G33), .B(new_n727_), .S(G29), .Z(new_n728_));
  XNOR2_X1  g303(.A(KEYINPUT57), .B(G2072), .ZN(new_n729_));
  XNOR2_X1  g304(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  NAND2_X1  g305(.A1(new_n684_), .A2(G27), .ZN(new_n731_));
  INV_X1    g306(.A(new_n494_), .ZN(new_n732_));
  OAI21_X1  g307(.A(new_n731_), .B1(new_n732_), .B2(new_n684_), .ZN(new_n733_));
  XOR2_X1   g308(.A(KEYINPUT68), .B(G2078), .Z(new_n734_));
  XNOR2_X1  g309(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NOR2_X1   g310(.A1(new_n730_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g311(.A1(new_n718_), .A2(new_n719_), .ZN(new_n737_));
  NOR2_X1   g312(.A1(G6), .A2(G16), .ZN(new_n738_));
  AOI21_X1  g313(.A(new_n738_), .B1(new_n557_), .B2(G16), .ZN(new_n739_));
  XOR2_X1   g314(.A(KEYINPUT70), .B(G1981), .Z(new_n740_));
  OR2_X1    g315(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g316(.A1(new_n739_), .A2(new_n740_), .ZN(new_n742_));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743_));
  OAI21_X1  g318(.A(G11), .B1(new_n743_), .B2(G868), .ZN(new_n744_));
  NOR2_X1   g319(.A1(KEYINPUT69), .A2(G28), .ZN(new_n745_));
  NOR2_X1   g320(.A1(new_n745_), .A2(G29), .ZN(new_n746_));
  NAND2_X1  g321(.A1(KEYINPUT69), .A2(G28), .ZN(new_n747_));
  AOI21_X1  g322(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g323(.A1(new_n737_), .A2(new_n741_), .A3(new_n742_), .A4(new_n748_), .ZN(new_n749_));
  AOI21_X1  g324(.A(new_n749_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n750_));
  NAND4_X1  g325(.A1(new_n699_), .A2(new_n721_), .A3(new_n736_), .A4(new_n750_), .ZN(new_n751_));
  NAND2_X1  g326(.A1(new_n709_), .A2(G1991), .ZN(new_n752_));
  AND3_X1   g327(.A1(new_n464_), .A2(new_n481_), .A3(G140), .ZN(new_n753_));
  XNOR2_X1  g328(.A(new_n753_), .B(KEYINPUT63), .ZN(new_n754_));
  AOI22_X1  g329(.A1(new_n464_), .A2(G128), .B1(G116), .B2(G2104), .ZN(new_n755_));
  NOR2_X1   g330(.A1(new_n755_), .A2(new_n471_), .ZN(new_n756_));
  NOR2_X1   g331(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g332(.A1(new_n482_), .A2(G104), .ZN(new_n758_));
  XOR2_X1   g333(.A(new_n758_), .B(KEYINPUT64), .Z(new_n759_));
  NAND2_X1  g334(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g335(.A1(new_n760_), .A2(G29), .ZN(new_n761_));
  NAND2_X1  g336(.A1(new_n684_), .A2(G26), .ZN(new_n762_));
  OR2_X1    g337(.A1(new_n762_), .A2(KEYINPUT62), .ZN(new_n763_));
  NAND2_X1  g338(.A1(new_n762_), .A2(KEYINPUT62), .ZN(new_n764_));
  NAND3_X1  g339(.A1(new_n761_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  XOR2_X1   g340(.A(KEYINPUT65), .B(G2067), .Z(new_n766_));
  OAI21_X1  g341(.A(new_n752_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g342(.A(new_n767_), .B1(new_n766_), .B2(new_n765_), .ZN(new_n768_));
  OR2_X1    g343(.A1(G29), .A2(G35), .ZN(new_n769_));
  OAI21_X1  g344(.A(new_n769_), .B1(new_n487_), .B2(new_n684_), .ZN(new_n770_));
  XNOR2_X1  g345(.A(KEYINPUT66), .B(G2090), .ZN(new_n771_));
  XNOR2_X1  g346(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  INV_X1    g347(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g348(.A(new_n768_), .B1(KEYINPUT67), .B2(new_n773_), .ZN(new_n774_));
  AOI211_X1 g349(.A(new_n751_), .B(new_n774_), .C1(KEYINPUT67), .C2(new_n773_), .ZN(new_n775_));
  INV_X1    g350(.A(KEYINPUT52), .ZN(new_n776_));
  OR2_X1    g351(.A1(new_n776_), .A2(G34), .ZN(new_n777_));
  NAND2_X1  g352(.A1(new_n776_), .A2(G34), .ZN(new_n778_));
  AOI21_X1  g353(.A(G29), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g354(.A(new_n779_), .B(KEYINPUT53), .ZN(new_n780_));
  INV_X1    g355(.A(KEYINPUT54), .ZN(new_n781_));
  OAI21_X1  g356(.A(new_n781_), .B1(new_n470_), .B2(new_n479_), .ZN(new_n782_));
  INV_X1    g357(.A(new_n476_), .ZN(new_n783_));
  AOI21_X1  g358(.A(new_n783_), .B1(new_n483_), .B2(G137), .ZN(new_n784_));
  NAND3_X1  g359(.A1(new_n467_), .A2(new_n468_), .A3(new_n465_), .ZN(new_n785_));
  NAND2_X1  g360(.A1(new_n785_), .A2(KEYINPUT10), .ZN(new_n786_));
  NAND3_X1  g361(.A1(new_n464_), .A2(new_n461_), .A3(new_n465_), .ZN(new_n787_));
  NAND2_X1  g362(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g363(.A1(new_n784_), .A2(KEYINPUT54), .A3(new_n788_), .A4(new_n475_), .ZN(new_n789_));
  NAND2_X1  g364(.A1(new_n782_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g365(.A(new_n780_), .B1(new_n790_), .B2(new_n684_), .ZN(new_n791_));
  XNOR2_X1  g366(.A(new_n791_), .B(KEYINPUT55), .ZN(new_n792_));
  INV_X1    g367(.A(G2084), .ZN(new_n793_));
  XNOR2_X1  g368(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  NAND2_X1  g369(.A1(new_n716_), .A2(G20), .ZN(new_n795_));
  XOR2_X1   g370(.A(new_n795_), .B(KEYINPUT48), .Z(new_n796_));
  OAI21_X1  g371(.A(new_n796_), .B1(new_n537_), .B2(new_n716_), .ZN(new_n797_));
  XNOR2_X1  g372(.A(new_n797_), .B(G1956), .ZN(new_n798_));
  NOR2_X1   g373(.A1(G5), .A2(G16), .ZN(new_n799_));
  AOI21_X1  g374(.A(new_n799_), .B1(G171), .B2(G16), .ZN(new_n800_));
  XNOR2_X1  g375(.A(new_n800_), .B(G1961), .ZN(new_n801_));
  NOR2_X1   g376(.A1(new_n798_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g377(.A1(new_n716_), .A2(G19), .ZN(new_n803_));
  XNOR2_X1  g378(.A(new_n803_), .B(KEYINPUT43), .ZN(new_n804_));
  AOI21_X1  g379(.A(new_n804_), .B1(new_n590_), .B2(G16), .ZN(new_n805_));
  XNOR2_X1  g380(.A(new_n805_), .B(KEYINPUT45), .ZN(new_n806_));
  XOR2_X1   g381(.A(KEYINPUT44), .B(G1341), .Z(new_n807_));
  INV_X1    g382(.A(new_n807_), .ZN(new_n808_));
  AND2_X1   g383(.A1(KEYINPUT46), .A2(G4), .ZN(new_n809_));
  NOR2_X1   g384(.A1(KEYINPUT46), .A2(G4), .ZN(new_n810_));
  OAI21_X1  g385(.A(new_n716_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g386(.A(new_n811_), .B1(new_n588_), .B2(new_n716_), .ZN(new_n812_));
  XOR2_X1   g387(.A(KEYINPUT47), .B(G1348), .Z(new_n813_));
  OAI221_X1 g388(.A(new_n802_), .B1(new_n806_), .B2(new_n808_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g389(.A1(KEYINPUT49), .A2(G21), .ZN(new_n815_));
  INV_X1    g390(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g391(.A1(KEYINPUT49), .A2(G21), .ZN(new_n817_));
  AOI21_X1  g392(.A(G16), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g393(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g394(.A(new_n819_), .B1(G168), .B2(new_n716_), .ZN(new_n820_));
  INV_X1    g395(.A(new_n820_), .ZN(new_n821_));
  XOR2_X1   g396(.A(KEYINPUT50), .B(G1966), .Z(new_n822_));
  AOI22_X1  g397(.A1(new_n821_), .A2(new_n822_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n823_));
  OAI21_X1  g398(.A(new_n823_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n824_));
  AOI211_X1 g399(.A(new_n814_), .B(new_n824_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n825_));
  XOR2_X1   g400(.A(new_n825_), .B(KEYINPUT51), .Z(new_n826_));
  NAND3_X1  g401(.A1(new_n775_), .A2(new_n794_), .A3(new_n826_), .ZN(G150));
  XNOR2_X1  g402(.A(G150), .B(KEYINPUT74), .ZN(G311));
  INV_X1    g403(.A(G67), .ZN(new_n829_));
  OAI21_X1  g404(.A(G651), .B1(new_n829_), .B2(G543), .ZN(new_n830_));
  NAND2_X1  g405(.A1(new_n502_), .A2(new_n496_), .ZN(new_n831_));
  OAI221_X1 g406(.A(new_n830_), .B1(G55), .B2(new_n502_), .C1(G93), .C2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g407(.A1(G80), .A2(G543), .A3(G651), .ZN(new_n833_));
  INV_X1    g408(.A(KEYINPUT75), .ZN(new_n834_));
  XNOR2_X1  g409(.A(new_n833_), .B(new_n834_), .ZN(new_n835_));
  NAND2_X1  g410(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g411(.A(new_n836_), .B1(KEYINPUT76), .B2(G860), .ZN(new_n837_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n838_));
  XNOR2_X1  g413(.A(new_n590_), .B(KEYINPUT77), .ZN(new_n839_));
  NOR3_X1   g414(.A1(new_n839_), .A2(new_n584_), .A3(new_n576_), .ZN(new_n840_));
  NOR2_X1   g415(.A1(new_n840_), .A2(G860), .ZN(new_n841_));
  OAI21_X1  g416(.A(new_n839_), .B1(new_n584_), .B2(new_n576_), .ZN(new_n842_));
  AOI21_X1  g417(.A(new_n838_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  MUX2_X1   g418(.A(new_n837_), .B(new_n836_), .S(new_n843_), .Z(G145));
  NAND2_X1  g419(.A1(new_n595_), .A2(G130), .ZN(new_n845_));
  XNOR2_X1  g420(.A(new_n845_), .B(KEYINPUT80), .ZN(new_n846_));
  AND3_X1   g421(.A1(G118), .A2(G2104), .A3(G2105), .ZN(new_n847_));
  NAND3_X1  g422(.A1(new_n482_), .A2(KEYINPUT79), .A3(G106), .ZN(new_n848_));
  INV_X1    g423(.A(KEYINPUT79), .ZN(new_n849_));
  INV_X1    g424(.A(G106), .ZN(new_n850_));
  OAI21_X1  g425(.A(new_n849_), .B1(new_n702_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g426(.A(new_n847_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n852_));
  AND3_X1   g427(.A1(new_n464_), .A2(new_n481_), .A3(G142), .ZN(new_n853_));
  INV_X1    g428(.A(KEYINPUT78), .ZN(new_n854_));
  XNOR2_X1  g429(.A(new_n853_), .B(new_n854_), .ZN(new_n855_));
  NAND3_X1  g430(.A1(new_n846_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g431(.A(new_n856_), .B(new_n727_), .ZN(new_n857_));
  NAND3_X1  g432(.A1(new_n784_), .A2(new_n788_), .A3(new_n475_), .ZN(new_n858_));
  XNOR2_X1  g433(.A(new_n857_), .B(new_n858_), .ZN(new_n859_));
  NAND3_X1  g434(.A1(new_n757_), .A2(new_n759_), .A3(new_n494_), .ZN(new_n860_));
  INV_X1    g435(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g436(.A(new_n494_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n862_));
  OAI21_X1  g437(.A(new_n695_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g438(.A1(new_n760_), .A2(new_n732_), .ZN(new_n864_));
  INV_X1    g439(.A(new_n695_), .ZN(new_n865_));
  NAND3_X1  g440(.A1(new_n864_), .A2(new_n865_), .A3(new_n860_), .ZN(new_n866_));
  XNOR2_X1  g441(.A(new_n708_), .B(KEYINPUT81), .ZN(new_n867_));
  NAND3_X1  g442(.A1(new_n863_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g443(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g444(.A(new_n867_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n870_));
  OAI21_X1  g445(.A(new_n859_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g446(.A(new_n487_), .B(new_n601_), .ZN(new_n872_));
  XOR2_X1   g447(.A(new_n605_), .B(KEYINPUT82), .Z(new_n873_));
  INV_X1    g448(.A(new_n873_), .ZN(new_n874_));
  XNOR2_X1  g449(.A(new_n872_), .B(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g450(.A(new_n857_), .B(G160), .ZN(new_n876_));
  INV_X1    g451(.A(new_n867_), .ZN(new_n877_));
  NOR3_X1   g452(.A1(new_n861_), .A2(new_n862_), .A3(new_n695_), .ZN(new_n878_));
  AOI21_X1  g453(.A(new_n865_), .B1(new_n864_), .B2(new_n860_), .ZN(new_n879_));
  OAI21_X1  g454(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g455(.A1(new_n876_), .A2(new_n868_), .A3(new_n880_), .ZN(new_n881_));
  NAND3_X1  g456(.A1(new_n871_), .A2(new_n875_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g457(.A(G37), .ZN(new_n883_));
  NAND2_X1  g458(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g459(.A(new_n875_), .B1(new_n871_), .B2(new_n881_), .ZN(new_n885_));
  NOR2_X1   g460(.A1(new_n884_), .A2(new_n885_), .ZN(G395));
  XNOR2_X1  g461(.A(new_n576_), .B(G299), .ZN(new_n887_));
  INV_X1    g462(.A(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g463(.A(new_n836_), .B(new_n590_), .ZN(new_n889_));
  NAND2_X1  g464(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g465(.A1(new_n890_), .A2(new_n589_), .ZN(new_n891_));
  XNOR2_X1  g466(.A(new_n891_), .B(KEYINPUT84), .ZN(new_n892_));
  NAND2_X1  g467(.A1(new_n887_), .A2(new_n889_), .ZN(new_n893_));
  XNOR2_X1  g468(.A(new_n889_), .B(KEYINPUT83), .ZN(new_n894_));
  OAI21_X1  g469(.A(new_n893_), .B1(new_n894_), .B2(new_n887_), .ZN(new_n895_));
  NAND2_X1  g470(.A1(new_n895_), .A2(new_n589_), .ZN(new_n896_));
  OR2_X1    g471(.A1(new_n894_), .A2(new_n888_), .ZN(new_n897_));
  OAI211_X1 g472(.A(new_n892_), .B(new_n896_), .C1(new_n589_), .C2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g473(.A(new_n898_), .B(KEYINPUT85), .ZN(new_n899_));
  XNOR2_X1  g474(.A(G288), .B(KEYINPUT87), .ZN(new_n900_));
  XNOR2_X1  g475(.A(new_n900_), .B(G290), .ZN(new_n901_));
  XNOR2_X1  g476(.A(new_n557_), .B(KEYINPUT86), .ZN(new_n902_));
  XNOR2_X1  g477(.A(G166), .B(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g478(.A(new_n901_), .B(new_n903_), .ZN(new_n904_));
  OR2_X1    g479(.A1(new_n899_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g480(.A(new_n581_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n906_));
  INV_X1    g481(.A(new_n836_), .ZN(new_n907_));
  AOI22_X1  g482(.A1(new_n905_), .A2(new_n906_), .B1(new_n581_), .B2(new_n907_), .ZN(G295));
  AOI22_X1  g483(.A1(new_n905_), .A2(new_n906_), .B1(new_n581_), .B2(new_n907_), .ZN(G331));
  INV_X1    g484(.A(new_n904_), .ZN(new_n910_));
  INV_X1    g485(.A(KEYINPUT89), .ZN(new_n911_));
  AND2_X1   g486(.A1(new_n895_), .A2(new_n911_), .ZN(new_n912_));
  XOR2_X1   g487(.A(G171), .B(KEYINPUT88), .Z(new_n913_));
  XNOR2_X1  g488(.A(new_n913_), .B(G168), .ZN(new_n914_));
  NAND3_X1  g489(.A1(new_n897_), .A2(new_n890_), .A3(new_n914_), .ZN(new_n915_));
  NOR2_X1   g490(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g491(.A(new_n914_), .B1(new_n895_), .B2(KEYINPUT89), .ZN(new_n917_));
  OAI21_X1  g492(.A(new_n910_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  AND2_X1   g493(.A1(new_n895_), .A2(KEYINPUT89), .ZN(new_n919_));
  OAI221_X1 g494(.A(new_n904_), .B1(new_n919_), .B2(new_n914_), .C1(new_n912_), .C2(new_n915_), .ZN(new_n920_));
  AND4_X1   g495(.A1(KEYINPUT90), .A2(new_n918_), .A3(new_n920_), .A4(new_n883_), .ZN(new_n921_));
  OAI22_X1  g496(.A1(new_n912_), .A2(new_n915_), .B1(new_n919_), .B2(new_n914_), .ZN(new_n922_));
  AOI21_X1  g497(.A(G37), .B1(new_n922_), .B2(new_n910_), .ZN(new_n923_));
  AOI21_X1  g498(.A(KEYINPUT90), .B1(new_n923_), .B2(new_n920_), .ZN(new_n924_));
  NOR2_X1   g499(.A1(new_n921_), .A2(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g500(.A(new_n925_), .B(KEYINPUT91), .ZN(G397));
  XNOR2_X1  g501(.A(KEYINPUT93), .B(G40), .ZN(new_n927_));
  AOI21_X1  g502(.A(new_n927_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n928_));
  XOR2_X1   g503(.A(KEYINPUT92), .B(G1384), .Z(new_n929_));
  NAND2_X1  g504(.A1(new_n494_), .A2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g505(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  OR2_X1    g506(.A1(new_n931_), .A2(KEYINPUT94), .ZN(new_n932_));
  INV_X1    g507(.A(KEYINPUT95), .ZN(new_n933_));
  AND2_X1   g508(.A1(new_n929_), .A2(G40), .ZN(new_n934_));
  NAND2_X1  g509(.A1(new_n494_), .A2(new_n934_), .ZN(new_n935_));
  OAI21_X1  g510(.A(new_n933_), .B1(new_n858_), .B2(new_n935_), .ZN(new_n936_));
  NAND4_X1  g511(.A1(G160), .A2(KEYINPUT95), .A3(new_n494_), .A4(new_n934_), .ZN(new_n937_));
  NAND2_X1  g512(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g513(.A1(new_n931_), .A2(KEYINPUT94), .ZN(new_n939_));
  AND3_X1   g514(.A1(new_n932_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  NOR2_X1   g515(.A1(new_n760_), .A2(G2067), .ZN(new_n941_));
  NAND2_X1  g516(.A1(new_n760_), .A2(G2067), .ZN(new_n942_));
  INV_X1    g517(.A(new_n942_), .ZN(new_n943_));
  OAI21_X1  g518(.A(new_n940_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g519(.A(KEYINPUT96), .ZN(new_n945_));
  XNOR2_X1  g520(.A(new_n944_), .B(new_n945_), .ZN(new_n946_));
  XOR2_X1   g521(.A(KEYINPUT97), .B(G1996), .Z(new_n947_));
  NAND3_X1  g522(.A1(new_n940_), .A2(new_n865_), .A3(new_n947_), .ZN(new_n948_));
  NOR2_X1   g523(.A1(new_n865_), .A2(new_n947_), .ZN(new_n949_));
  NAND2_X1  g524(.A1(new_n940_), .A2(new_n949_), .ZN(new_n950_));
  INV_X1    g525(.A(KEYINPUT98), .ZN(new_n951_));
  AND3_X1   g526(.A1(new_n948_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  AOI21_X1  g527(.A(new_n951_), .B1(new_n948_), .B2(new_n950_), .ZN(new_n953_));
  NOR2_X1   g528(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  INV_X1    g529(.A(new_n940_), .ZN(new_n955_));
  NOR3_X1   g530(.A1(new_n955_), .A2(G1991), .A3(new_n708_), .ZN(new_n956_));
  AND2_X1   g531(.A1(new_n954_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g532(.A(new_n948_), .ZN(new_n958_));
  OAI21_X1  g533(.A(new_n946_), .B1(new_n957_), .B2(new_n958_), .ZN(new_n959_));
  XNOR2_X1  g534(.A(new_n708_), .B(G1991), .ZN(new_n960_));
  NAND2_X1  g535(.A1(new_n940_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g536(.A1(G290), .A2(G1986), .ZN(new_n962_));
  NAND2_X1  g537(.A1(new_n940_), .A2(new_n962_), .ZN(new_n963_));
  INV_X1    g538(.A(new_n963_), .ZN(new_n964_));
  NAND4_X1  g539(.A1(new_n954_), .A2(new_n946_), .A3(new_n961_), .A4(new_n964_), .ZN(new_n965_));
  NAND2_X1  g540(.A1(new_n940_), .A2(new_n941_), .ZN(new_n966_));
  XOR2_X1   g541(.A(new_n966_), .B(KEYINPUT99), .Z(new_n967_));
  NAND4_X1  g542(.A1(new_n959_), .A2(KEYINPUT100), .A3(new_n965_), .A4(new_n967_), .ZN(new_n968_));
  AOI21_X1  g543(.A(new_n958_), .B1(new_n954_), .B2(new_n956_), .ZN(new_n969_));
  INV_X1    g544(.A(new_n946_), .ZN(new_n970_));
  OAI211_X1 g545(.A(new_n965_), .B(new_n967_), .C1(new_n969_), .C2(new_n970_), .ZN(new_n971_));
  INV_X1    g546(.A(KEYINPUT100), .ZN(new_n972_));
  NAND2_X1  g547(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g548(.A1(new_n968_), .A2(new_n973_), .ZN(new_n974_));
  NAND2_X1  g549(.A1(G290), .A2(G1986), .ZN(new_n975_));
  INV_X1    g550(.A(new_n975_), .ZN(new_n976_));
  OAI21_X1  g551(.A(new_n940_), .B1(new_n962_), .B2(new_n976_), .ZN(new_n977_));
  INV_X1    g552(.A(KEYINPUT123), .ZN(new_n978_));
  XNOR2_X1  g553(.A(new_n977_), .B(new_n978_), .ZN(new_n979_));
  NAND4_X1  g554(.A1(new_n954_), .A2(new_n946_), .A3(new_n979_), .A4(new_n961_), .ZN(new_n980_));
  XNOR2_X1  g555(.A(new_n980_), .B(KEYINPUT124), .ZN(new_n981_));
  INV_X1    g556(.A(G1981), .ZN(new_n982_));
  NAND4_X1  g557(.A1(new_n938_), .A2(G8), .A3(new_n982_), .A4(G305), .ZN(new_n983_));
  XNOR2_X1  g558(.A(new_n983_), .B(KEYINPUT101), .ZN(new_n984_));
  INV_X1    g559(.A(G8), .ZN(new_n985_));
  AOI21_X1  g560(.A(new_n985_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n986_));
  OAI21_X1  g561(.A(new_n986_), .B1(new_n982_), .B2(G305), .ZN(new_n987_));
  INV_X1    g562(.A(new_n987_), .ZN(new_n988_));
  NAND2_X1  g563(.A1(new_n984_), .A2(new_n988_), .ZN(new_n989_));
  XOR2_X1   g564(.A(KEYINPUT106), .B(G1976), .Z(new_n990_));
  AND2_X1   g565(.A1(new_n986_), .A2(new_n990_), .ZN(new_n991_));
  NAND2_X1  g566(.A1(new_n938_), .A2(G288), .ZN(new_n992_));
  NAND2_X1  g567(.A1(new_n992_), .A2(KEYINPUT121), .ZN(new_n993_));
  OR2_X1    g568(.A1(new_n992_), .A2(KEYINPUT121), .ZN(new_n994_));
  NAND4_X1  g569(.A1(new_n989_), .A2(new_n991_), .A3(new_n993_), .A4(new_n994_), .ZN(new_n995_));
  NAND4_X1  g570(.A1(new_n938_), .A2(G8), .A3(G288), .A4(new_n990_), .ZN(new_n996_));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n997_));
  NAND2_X1  g572(.A1(new_n996_), .A2(new_n997_), .ZN(new_n998_));
  NAND4_X1  g573(.A1(new_n986_), .A2(KEYINPUT107), .A3(G288), .A4(new_n990_), .ZN(new_n999_));
  NAND2_X1  g574(.A1(new_n938_), .A2(G8), .ZN(new_n1000_));
  NOR2_X1   g575(.A1(G288), .A2(new_n990_), .ZN(new_n1001_));
  NOR2_X1   g576(.A1(new_n1000_), .A2(new_n1001_), .ZN(new_n1002_));
  NAND3_X1  g577(.A1(new_n998_), .A2(new_n999_), .A3(new_n1002_), .ZN(new_n1003_));
  NAND2_X1  g578(.A1(new_n1003_), .A2(KEYINPUT108), .ZN(new_n1004_));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n1005_));
  NAND4_X1  g580(.A1(new_n998_), .A2(new_n1002_), .A3(new_n1005_), .A4(new_n999_), .ZN(new_n1006_));
  NAND2_X1  g581(.A1(new_n1004_), .A2(new_n1006_), .ZN(new_n1007_));
  XNOR2_X1  g582(.A(KEYINPUT110), .B(G1961), .ZN(new_n1008_));
  INV_X1    g583(.A(new_n1008_), .ZN(new_n1009_));
  NAND3_X1  g584(.A1(new_n494_), .A2(KEYINPUT102), .A3(new_n929_), .ZN(new_n1010_));
  NAND3_X1  g585(.A1(new_n1010_), .A2(G160), .A3(G40), .ZN(new_n1011_));
  INV_X1    g586(.A(new_n1011_), .ZN(new_n1012_));
  AOI21_X1  g587(.A(KEYINPUT102), .B1(new_n494_), .B2(new_n929_), .ZN(new_n1013_));
  INV_X1    g588(.A(new_n1013_), .ZN(new_n1014_));
  AOI21_X1  g589(.A(new_n1009_), .B1(new_n1012_), .B2(new_n1014_), .ZN(new_n1015_));
  INV_X1    g590(.A(G2078), .ZN(new_n1016_));
  INV_X1    g591(.A(new_n930_), .ZN(new_n1017_));
  INV_X1    g592(.A(new_n927_), .ZN(new_n1018_));
  NAND4_X1  g593(.A1(new_n790_), .A2(new_n1016_), .A3(new_n1017_), .A4(new_n1018_), .ZN(new_n1019_));
  NAND2_X1  g594(.A1(new_n1019_), .A2(KEYINPUT109), .ZN(new_n1020_));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n1021_));
  NAND4_X1  g596(.A1(new_n928_), .A2(new_n1021_), .A3(new_n1016_), .A4(new_n1017_), .ZN(new_n1022_));
  AOI211_X1 g597(.A(G171), .B(new_n1015_), .C1(new_n1020_), .C2(new_n1022_), .ZN(new_n1023_));
  NAND2_X1  g598(.A1(new_n1020_), .A2(new_n1022_), .ZN(new_n1024_));
  INV_X1    g599(.A(new_n1015_), .ZN(new_n1025_));
  AOI21_X1  g600(.A(G301), .B1(new_n1024_), .B2(new_n1025_), .ZN(new_n1026_));
  OAI21_X1  g601(.A(KEYINPUT111), .B1(new_n1023_), .B2(new_n1026_), .ZN(new_n1027_));
  NAND2_X1  g602(.A1(new_n1024_), .A2(new_n1025_), .ZN(new_n1028_));
  NAND2_X1  g603(.A1(new_n1028_), .A2(G171), .ZN(new_n1029_));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n1030_));
  NAND3_X1  g605(.A1(new_n1024_), .A2(G301), .A3(new_n1025_), .ZN(new_n1031_));
  NAND3_X1  g606(.A1(new_n1029_), .A2(new_n1030_), .A3(new_n1031_), .ZN(new_n1032_));
  AND3_X1   g607(.A1(new_n1007_), .A2(new_n1027_), .A3(new_n1032_), .ZN(new_n1033_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n1034_));
  INV_X1    g609(.A(G1956), .ZN(new_n1035_));
  OAI21_X1  g610(.A(new_n1035_), .B1(new_n1011_), .B2(new_n1013_), .ZN(new_n1036_));
  INV_X1    g611(.A(G2072), .ZN(new_n1037_));
  NAND4_X1  g612(.A1(new_n790_), .A2(new_n1037_), .A3(new_n1017_), .A4(new_n1018_), .ZN(new_n1038_));
  NAND2_X1  g613(.A1(new_n1036_), .A2(new_n1038_), .ZN(new_n1039_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n1040_));
  AOI21_X1  g615(.A(G299), .B1(new_n1039_), .B2(new_n1040_), .ZN(new_n1041_));
  NAND3_X1  g616(.A1(new_n1036_), .A2(new_n1038_), .A3(KEYINPUT115), .ZN(new_n1042_));
  AND3_X1   g617(.A1(new_n1041_), .A2(KEYINPUT116), .A3(new_n1042_), .ZN(new_n1043_));
  AOI21_X1  g618(.A(KEYINPUT116), .B1(new_n1041_), .B2(new_n1042_), .ZN(new_n1044_));
  NOR2_X1   g619(.A1(new_n1043_), .A2(new_n1044_), .ZN(new_n1045_));
  NAND2_X1  g620(.A1(new_n1039_), .A2(new_n537_), .ZN(new_n1046_));
  NAND3_X1  g621(.A1(new_n1036_), .A2(new_n1038_), .A3(G299), .ZN(new_n1047_));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048_));
  INV_X1    g623(.A(G1348), .ZN(new_n1049_));
  OAI21_X1  g624(.A(new_n1049_), .B1(new_n1011_), .B2(new_n1013_), .ZN(new_n1050_));
  INV_X1    g625(.A(G2067), .ZN(new_n1051_));
  NAND4_X1  g626(.A1(new_n790_), .A2(new_n1051_), .A3(new_n1017_), .A4(new_n1018_), .ZN(new_n1052_));
  AOI21_X1  g627(.A(new_n576_), .B1(new_n1050_), .B2(new_n1052_), .ZN(new_n1053_));
  OAI211_X1 g628(.A(new_n1046_), .B(new_n1047_), .C1(new_n1048_), .C2(new_n1053_), .ZN(new_n1054_));
  NAND2_X1  g629(.A1(new_n1053_), .A2(new_n1048_), .ZN(new_n1055_));
  INV_X1    g630(.A(new_n1055_), .ZN(new_n1056_));
  XOR2_X1   g631(.A(KEYINPUT117), .B(G1341), .Z(new_n1057_));
  NAND2_X1  g632(.A1(new_n938_), .A2(new_n1057_), .ZN(new_n1058_));
  NAND3_X1  g633(.A1(new_n928_), .A2(new_n1017_), .A3(new_n947_), .ZN(new_n1059_));
  AOI21_X1  g634(.A(new_n590_), .B1(new_n1058_), .B2(new_n1059_), .ZN(new_n1060_));
  NAND3_X1  g635(.A1(new_n1060_), .A2(new_n1046_), .A3(new_n1047_), .ZN(new_n1061_));
  AND3_X1   g636(.A1(new_n1050_), .A2(new_n1052_), .A3(new_n577_), .ZN(new_n1062_));
  AOI21_X1  g637(.A(new_n577_), .B1(new_n1050_), .B2(new_n1052_), .ZN(new_n1063_));
  NOR2_X1   g638(.A1(new_n1062_), .A2(new_n1063_), .ZN(new_n1064_));
  OAI22_X1  g639(.A1(new_n1054_), .A2(new_n1056_), .B1(new_n1061_), .B2(new_n1064_), .ZN(new_n1065_));
  OAI21_X1  g640(.A(new_n1034_), .B1(new_n1045_), .B2(new_n1065_), .ZN(new_n1066_));
  NAND2_X1  g641(.A1(new_n1041_), .A2(new_n1042_), .ZN(new_n1067_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068_));
  NAND2_X1  g643(.A1(new_n1067_), .A2(new_n1068_), .ZN(new_n1069_));
  NAND3_X1  g644(.A1(new_n1041_), .A2(KEYINPUT116), .A3(new_n1042_), .ZN(new_n1070_));
  NAND2_X1  g645(.A1(new_n1069_), .A2(new_n1070_), .ZN(new_n1071_));
  OR2_X1    g646(.A1(new_n1061_), .A2(new_n1064_), .ZN(new_n1072_));
  OR2_X1    g647(.A1(new_n1053_), .A2(new_n1048_), .ZN(new_n1073_));
  NAND4_X1  g648(.A1(new_n1073_), .A2(new_n1046_), .A3(new_n1047_), .A4(new_n1055_), .ZN(new_n1074_));
  NAND4_X1  g649(.A1(new_n1071_), .A2(KEYINPUT118), .A3(new_n1072_), .A4(new_n1074_), .ZN(new_n1075_));
  NAND3_X1  g650(.A1(new_n1033_), .A2(new_n1066_), .A3(new_n1075_), .ZN(new_n1076_));
  INV_X1    g651(.A(KEYINPUT103), .ZN(new_n1077_));
  NAND4_X1  g652(.A1(new_n1014_), .A2(G40), .A3(G160), .A4(new_n1010_), .ZN(new_n1078_));
  OAI21_X1  g653(.A(new_n1077_), .B1(new_n1078_), .B2(G2084), .ZN(new_n1079_));
  NAND4_X1  g654(.A1(new_n1012_), .A2(KEYINPUT103), .A3(new_n793_), .A4(new_n1014_), .ZN(new_n1080_));
  NAND3_X1  g655(.A1(new_n790_), .A2(new_n1017_), .A3(new_n1018_), .ZN(new_n1081_));
  INV_X1    g656(.A(G1966), .ZN(new_n1082_));
  NAND2_X1  g657(.A1(new_n1081_), .A2(new_n1082_), .ZN(new_n1083_));
  NAND3_X1  g658(.A1(new_n1079_), .A2(new_n1080_), .A3(new_n1083_), .ZN(new_n1084_));
  NAND2_X1  g659(.A1(new_n1084_), .A2(G8), .ZN(new_n1085_));
  NAND2_X1  g660(.A1(G286), .A2(G8), .ZN(new_n1086_));
  XNOR2_X1  g661(.A(new_n1086_), .B(KEYINPUT104), .ZN(new_n1087_));
  INV_X1    g662(.A(new_n1087_), .ZN(new_n1088_));
  NAND2_X1  g663(.A1(new_n1085_), .A2(new_n1088_), .ZN(new_n1089_));
  NAND3_X1  g664(.A1(new_n1084_), .A2(new_n1087_), .A3(G8), .ZN(new_n1090_));
  NAND3_X1  g665(.A1(new_n989_), .A2(new_n1089_), .A3(new_n1090_), .ZN(new_n1091_));
  NAND2_X1  g666(.A1(new_n1091_), .A2(KEYINPUT105), .ZN(new_n1092_));
  NAND2_X1  g667(.A1(G303), .A2(G8), .ZN(new_n1093_));
  NOR2_X1   g668(.A1(new_n1078_), .A2(G2090), .ZN(new_n1094_));
  AOI21_X1  g669(.A(G1971), .B1(new_n928_), .B2(new_n1017_), .ZN(new_n1095_));
  OAI21_X1  g670(.A(G8), .B1(new_n1094_), .B2(new_n1095_), .ZN(new_n1096_));
  INV_X1    g671(.A(G1971), .ZN(new_n1097_));
  NAND2_X1  g672(.A1(new_n1081_), .A2(new_n1097_), .ZN(new_n1098_));
  INV_X1    g673(.A(G2090), .ZN(new_n1099_));
  NAND3_X1  g674(.A1(new_n1012_), .A2(new_n1099_), .A3(new_n1014_), .ZN(new_n1100_));
  AOI21_X1  g675(.A(new_n1093_), .B1(new_n1098_), .B2(new_n1100_), .ZN(new_n1101_));
  AOI22_X1  g676(.A1(new_n1093_), .A2(new_n1096_), .B1(new_n1101_), .B2(KEYINPUT112), .ZN(new_n1102_));
  NOR2_X1   g677(.A1(new_n1101_), .A2(KEYINPUT112), .ZN(new_n1103_));
  INV_X1    g678(.A(new_n1103_), .ZN(new_n1104_));
  NAND3_X1  g679(.A1(new_n1102_), .A2(new_n1104_), .A3(KEYINPUT113), .ZN(new_n1105_));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n1106_));
  INV_X1    g681(.A(new_n1093_), .ZN(new_n1107_));
  OAI211_X1 g682(.A(KEYINPUT112), .B(new_n1107_), .C1(new_n1094_), .C2(new_n1095_), .ZN(new_n1108_));
  AOI21_X1  g683(.A(new_n985_), .B1(new_n1098_), .B2(new_n1100_), .ZN(new_n1109_));
  OAI21_X1  g684(.A(new_n1108_), .B1(new_n1107_), .B2(new_n1109_), .ZN(new_n1110_));
  OAI21_X1  g685(.A(new_n1106_), .B1(new_n1110_), .B2(new_n1103_), .ZN(new_n1111_));
  NAND2_X1  g686(.A1(new_n1105_), .A2(new_n1111_), .ZN(new_n1112_));
  INV_X1    g687(.A(KEYINPUT105), .ZN(new_n1113_));
  NAND4_X1  g688(.A1(new_n989_), .A2(new_n1113_), .A3(new_n1089_), .A4(new_n1090_), .ZN(new_n1114_));
  NAND3_X1  g689(.A1(new_n1092_), .A2(new_n1112_), .A3(new_n1114_), .ZN(new_n1115_));
  OAI21_X1  g690(.A(new_n995_), .B1(new_n1076_), .B2(new_n1115_), .ZN(new_n1116_));
  INV_X1    g691(.A(new_n1090_), .ZN(new_n1117_));
  OR2_X1    g692(.A1(new_n983_), .A2(KEYINPUT101), .ZN(new_n1118_));
  NAND2_X1  g693(.A1(new_n983_), .A2(KEYINPUT101), .ZN(new_n1119_));
  AOI21_X1  g694(.A(new_n987_), .B1(new_n1118_), .B2(new_n1119_), .ZN(new_n1120_));
  AOI21_X1  g695(.A(new_n1087_), .B1(new_n1084_), .B2(G8), .ZN(new_n1121_));
  NOR3_X1   g696(.A1(new_n1117_), .A2(new_n1120_), .A3(new_n1121_), .ZN(new_n1122_));
  NOR2_X1   g697(.A1(new_n1029_), .A2(KEYINPUT119), .ZN(new_n1123_));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124_));
  OAI21_X1  g699(.A(new_n1003_), .B1(new_n1026_), .B2(new_n1124_), .ZN(new_n1125_));
  NOR2_X1   g700(.A1(new_n1123_), .A2(new_n1125_), .ZN(new_n1126_));
  NAND3_X1  g701(.A1(new_n1112_), .A2(new_n1122_), .A3(new_n1126_), .ZN(new_n1127_));
  NOR2_X1   g702(.A1(new_n1120_), .A2(new_n1090_), .ZN(new_n1128_));
  NAND3_X1  g703(.A1(new_n1112_), .A2(new_n1007_), .A3(new_n1128_), .ZN(new_n1129_));
  NOR3_X1   g704(.A1(new_n1000_), .A2(G1981), .A3(G305), .ZN(new_n1130_));
  NOR3_X1   g705(.A1(new_n1120_), .A2(G303), .A3(new_n1096_), .ZN(new_n1131_));
  AOI21_X1  g706(.A(new_n1130_), .B1(new_n1131_), .B2(new_n1007_), .ZN(new_n1132_));
  NAND3_X1  g707(.A1(new_n1127_), .A2(new_n1129_), .A3(new_n1132_), .ZN(new_n1133_));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n1134_));
  NAND2_X1  g709(.A1(new_n1133_), .A2(new_n1134_), .ZN(new_n1135_));
  NAND4_X1  g710(.A1(new_n1127_), .A2(new_n1129_), .A3(KEYINPUT120), .A4(new_n1132_), .ZN(new_n1136_));
  AOI21_X1  g711(.A(new_n1116_), .B1(new_n1135_), .B2(new_n1136_), .ZN(new_n1137_));
  OAI21_X1  g712(.A(new_n981_), .B1(new_n1137_), .B2(KEYINPUT122), .ZN(new_n1138_));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139_));
  AOI211_X1 g714(.A(new_n1139_), .B(new_n1116_), .C1(new_n1135_), .C2(new_n1136_), .ZN(new_n1140_));
  OAI21_X1  g715(.A(new_n974_), .B1(new_n1138_), .B2(new_n1140_), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g716(.A(new_n650_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n1143_));
  NAND2_X1  g717(.A1(new_n1143_), .A2(KEYINPUT125), .ZN(new_n1144_));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1145_));
  OAI211_X1 g719(.A(new_n1145_), .B(new_n650_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n1146_));
  NAND2_X1  g720(.A1(new_n1144_), .A2(new_n1146_), .ZN(new_n1147_));
  OAI21_X1  g721(.A(new_n633_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n1148_));
  NAND2_X1  g722(.A1(new_n1148_), .A2(KEYINPUT126), .ZN(new_n1149_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1150_));
  OAI211_X1 g724(.A(new_n633_), .B(new_n1150_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n1151_));
  NAND3_X1  g725(.A1(new_n1149_), .A2(G319), .A3(new_n1151_), .ZN(new_n1152_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n1152_), .ZN(new_n1153_));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1154_));
  AND3_X1   g728(.A1(new_n1147_), .A2(new_n1153_), .A3(new_n1154_), .ZN(new_n1155_));
  AOI21_X1  g729(.A(new_n1154_), .B1(new_n1147_), .B2(new_n1153_), .ZN(new_n1156_));
  NOR2_X1   g730(.A1(new_n1155_), .A2(new_n1156_), .ZN(G308));
  NAND2_X1  g731(.A1(new_n1147_), .A2(new_n1153_), .ZN(G225));
endmodule


