//Secret key is'1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_c6288" written by ABC on Wed Nov 16 10:20:01 2022

module locked_c6288 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1gat, G18gat, G35gat, G52gat, G69gat,
    G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat,
    G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat,
    G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat,
    G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1gat, G18gat, G35gat, G52gat,
    G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat,
    G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat,
    G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat,
    G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_n193_, new_n194_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_,
    new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_,
    new_n2725_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2907_, new_n2908_;
  INV_X1    g0000(.A(G1gat), .ZN(new_n193_));
  INV_X1    g0001(.A(G273gat), .ZN(new_n194_));
  NOR2_X1   g0002(.A1(new_n193_), .A2(new_n194_), .ZN(G545gat));
  INV_X1    g0003(.A(G18gat), .ZN(new_n196_));
  NOR2_X1   g0004(.A1(new_n196_), .A2(new_n194_), .ZN(new_n197_));
  INV_X1    g0005(.A(G290gat), .ZN(new_n198_));
  NOR2_X1   g0006(.A1(new_n193_), .A2(new_n198_), .ZN(new_n199_));
  XOR2_X1   g0007(.A(new_n197_), .B(new_n199_), .Z(G1581gat));
  NAND3_X1  g0008(.A1(new_n197_), .A2(G35gat), .A3(G290gat), .ZN(new_n201_));
  NAND2_X1  g0009(.A1(new_n201_), .A2(KEYINPUT0), .ZN(new_n202_));
  AOI22_X1  g0010(.A1(G18gat), .A2(G290gat), .B1(G35gat), .B2(G273gat), .ZN(new_n203_));
  AND2_X1   g0011(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g0012(.A1(new_n197_), .A2(new_n199_), .ZN(new_n205_));
  OAI21_X1  g0013(.A(new_n205_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n206_));
  NOR2_X1   g0014(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g0015(.A1(new_n202_), .A2(new_n205_), .ZN(new_n208_));
  NOR2_X1   g0016(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g0017(.A1(G1gat), .A2(G307gat), .ZN(new_n210_));
  XNOR2_X1  g0018(.A(new_n209_), .B(new_n210_), .ZN(G1901gat));
  INV_X1    g0019(.A(new_n201_), .ZN(new_n212_));
  INV_X1    g0020(.A(G35gat), .ZN(new_n213_));
  INV_X1    g0021(.A(G52gat), .ZN(new_n214_));
  OAI22_X1  g0022(.A1(new_n213_), .A2(new_n198_), .B1(new_n214_), .B2(new_n194_), .ZN(new_n215_));
  NAND4_X1  g0023(.A1(G35gat), .A2(G52gat), .A3(G273gat), .A4(G290gat), .ZN(new_n216_));
  NAND2_X1  g0024(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g0025(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n218_));
  INV_X1    g0026(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g0027(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n220_));
  AOI21_X1  g0028(.A(new_n212_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g0029(.A1(new_n218_), .A2(new_n201_), .ZN(new_n222_));
  NOR2_X1   g0030(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g0031(.A1(G18gat), .A2(G307gat), .ZN(new_n224_));
  XNOR2_X1  g0032(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g0033(.A1(new_n209_), .A2(new_n210_), .ZN(new_n226_));
  OAI21_X1  g0034(.A(new_n226_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n227_));
  NAND2_X1  g0035(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g0036(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g0037(.A1(new_n225_), .A2(new_n227_), .ZN(new_n230_));
  NOR2_X1   g0038(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g0039(.A(G324gat), .ZN(new_n232_));
  NOR2_X1   g0040(.A1(new_n193_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g0041(.A(new_n231_), .B(new_n233_), .Z(G2223gat));
  OAI21_X1  g0042(.A(new_n224_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n235_));
  NAND2_X1  g0043(.A1(new_n217_), .A2(new_n201_), .ZN(new_n236_));
  XNOR2_X1  g0044(.A(new_n236_), .B(KEYINPUT2), .ZN(new_n237_));
  NAND2_X1  g0045(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g0046(.A1(G52gat), .A2(G69gat), .A3(G273gat), .A4(G290gat), .ZN(new_n239_));
  INV_X1    g0047(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g0048(.A1(new_n240_), .A2(new_n216_), .ZN(new_n241_));
  AOI22_X1  g0049(.A1(G52gat), .A2(G290gat), .B1(G69gat), .B2(G273gat), .ZN(new_n242_));
  OR2_X1    g0050(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g0051(.A(new_n241_), .B1(new_n243_), .B2(new_n216_), .ZN(new_n244_));
  INV_X1    g0052(.A(G307gat), .ZN(new_n245_));
  NOR2_X1   g0053(.A1(new_n213_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g0054(.A(new_n244_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g0055(.A1(new_n238_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g0056(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g0057(.A1(new_n238_), .A2(new_n247_), .ZN(new_n250_));
  NOR2_X1   g0058(.A1(new_n196_), .A2(new_n232_), .ZN(new_n251_));
  OR3_X1    g0059(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g0060(.A(new_n251_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n253_));
  NAND2_X1  g0061(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g0062(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g0063(.A(new_n228_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n256_));
  NAND2_X1  g0064(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g0065(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g0066(.A1(new_n255_), .A2(new_n256_), .ZN(new_n259_));
  NOR2_X1   g0067(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g0068(.A(G341gat), .ZN(new_n261_));
  NOR2_X1   g0069(.A1(new_n193_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g0070(.A(new_n260_), .B(new_n262_), .Z(G2548gat));
  NAND2_X1  g0071(.A1(new_n252_), .A2(new_n248_), .ZN(new_n264_));
  NAND4_X1  g0072(.A1(G69gat), .A2(G86gat), .A3(G273gat), .A4(G290gat), .ZN(new_n265_));
  INV_X1    g0073(.A(new_n265_), .ZN(new_n266_));
  AOI22_X1  g0074(.A1(G69gat), .A2(G290gat), .B1(G86gat), .B2(G273gat), .ZN(new_n267_));
  OAI21_X1  g0075(.A(new_n239_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g0076(.A1(new_n240_), .A2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g0077(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g0078(.A1(G52gat), .A2(G307gat), .ZN(new_n271_));
  XNOR2_X1  g0079(.A(new_n271_), .B(KEYINPUT3), .ZN(new_n272_));
  XNOR2_X1  g0080(.A(new_n270_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g0081(.A1(new_n243_), .A2(new_n216_), .ZN(new_n274_));
  OAI21_X1  g0082(.A(new_n274_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n275_));
  NOR2_X1   g0083(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g0084(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g0085(.A1(new_n273_), .A2(new_n275_), .ZN(new_n278_));
  NAND2_X1  g0086(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g0087(.A1(new_n213_), .A2(new_n232_), .ZN(new_n280_));
  INV_X1    g0088(.A(KEYINPUT4), .ZN(new_n281_));
  XNOR2_X1  g0089(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  NAND2_X1  g0090(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  OAI211_X1 g0091(.A(new_n277_), .B(new_n278_), .C1(new_n281_), .C2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g0092(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g0093(.A1(new_n264_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g0094(.A1(G18gat), .A2(G341gat), .ZN(new_n287_));
  NAND4_X1  g0095(.A1(new_n252_), .A2(new_n248_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n288_));
  NAND3_X1  g0096(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g0097(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g0098(.A(new_n287_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n291_));
  NOR2_X1   g0099(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g0100(.A(new_n257_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n293_));
  NOR2_X1   g0101(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g0102(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g0103(.A1(new_n292_), .A2(new_n293_), .ZN(new_n296_));
  NAND2_X1  g0104(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g0105(.A(KEYINPUT5), .ZN(new_n298_));
  NAND2_X1  g0106(.A1(new_n298_), .A2(G358gat), .ZN(new_n299_));
  INV_X1    g0107(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g0108(.A1(new_n298_), .A2(G358gat), .ZN(new_n301_));
  NOR2_X1   g0109(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g0110(.A1(new_n302_), .A2(new_n193_), .ZN(new_n303_));
  XNOR2_X1  g0111(.A(new_n297_), .B(new_n303_), .ZN(G2877gat));
  OAI21_X1  g0112(.A(new_n296_), .B1(new_n294_), .B2(new_n303_), .ZN(new_n305_));
  AOI21_X1  g0113(.A(new_n276_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n306_));
  INV_X1    g0114(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g0115(.A1(G103gat), .A2(G290gat), .ZN(new_n308_));
  INV_X1    g0116(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g0117(.A1(new_n309_), .A2(G86gat), .A3(G273gat), .ZN(new_n310_));
  NAND2_X1  g0118(.A1(G103gat), .A2(G273gat), .ZN(new_n311_));
  INV_X1    g0119(.A(G86gat), .ZN(new_n312_));
  OAI21_X1  g0120(.A(new_n311_), .B1(new_n312_), .B2(new_n198_), .ZN(new_n313_));
  NAND2_X1  g0121(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g0122(.A1(new_n314_), .A2(new_n265_), .ZN(new_n315_));
  NAND2_X1  g0123(.A1(new_n310_), .A2(new_n266_), .ZN(new_n316_));
  NAND2_X1  g0124(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g0125(.A(G69gat), .ZN(new_n318_));
  NOR2_X1   g0126(.A1(new_n318_), .A2(new_n245_), .ZN(new_n319_));
  NAND2_X1  g0127(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g0128(.A1(new_n268_), .A2(new_n272_), .A3(new_n269_), .ZN(new_n321_));
  NAND2_X1  g0129(.A1(new_n321_), .A2(new_n268_), .ZN(new_n322_));
  INV_X1    g0130(.A(new_n319_), .ZN(new_n323_));
  NAND3_X1  g0131(.A1(new_n315_), .A2(new_n316_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g0132(.A1(new_n320_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g0133(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g0134(.A(new_n322_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n327_));
  NOR2_X1   g0135(.A1(new_n214_), .A2(new_n232_), .ZN(new_n328_));
  NOR3_X1   g0136(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g0137(.A(new_n328_), .ZN(new_n330_));
  INV_X1    g0138(.A(new_n327_), .ZN(new_n331_));
  AOI21_X1  g0139(.A(new_n330_), .B1(new_n331_), .B2(new_n325_), .ZN(new_n332_));
  NOR3_X1   g0140(.A1(new_n307_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g0141(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g0142(.A1(new_n213_), .A2(new_n261_), .ZN(new_n335_));
  INV_X1    g0143(.A(new_n335_), .ZN(new_n336_));
  OAI21_X1  g0144(.A(new_n307_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n337_));
  NAND3_X1  g0145(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g0146(.A(new_n337_), .ZN(new_n339_));
  OAI21_X1  g0147(.A(new_n335_), .B1(new_n339_), .B2(new_n333_), .ZN(new_n340_));
  AND2_X1   g0148(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g0149(.A1(new_n289_), .A2(KEYINPUT6), .ZN(new_n342_));
  INV_X1    g0150(.A(new_n286_), .ZN(new_n343_));
  AOI21_X1  g0151(.A(new_n343_), .B1(new_n289_), .B2(KEYINPUT6), .ZN(new_n344_));
  AOI21_X1  g0152(.A(new_n341_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g0153(.A1(new_n289_), .A2(new_n286_), .A3(new_n341_), .ZN(new_n346_));
  INV_X1    g0154(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g0155(.A(new_n302_), .ZN(new_n348_));
  NAND2_X1  g0156(.A1(new_n348_), .A2(G18gat), .ZN(new_n349_));
  OR3_X1    g0157(.A1(new_n345_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  OAI21_X1  g0158(.A(new_n349_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n351_));
  AOI21_X1  g0159(.A(new_n305_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g0160(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g0161(.A1(new_n350_), .A2(new_n305_), .A3(new_n351_), .ZN(new_n354_));
  NAND2_X1  g0162(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g0163(.A(G375gat), .ZN(new_n356_));
  NOR2_X1   g0164(.A1(new_n193_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g0165(.A(new_n355_), .B(new_n357_), .ZN(G3211gat));
  NOR2_X1   g0166(.A1(new_n196_), .A2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g0167(.A1(new_n342_), .A2(new_n344_), .ZN(new_n360_));
  NAND2_X1  g0168(.A1(new_n360_), .A2(new_n341_), .ZN(new_n361_));
  NOR2_X1   g0169(.A1(new_n302_), .A2(new_n213_), .ZN(new_n362_));
  AOI21_X1  g0170(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n363_));
  OAI21_X1  g0171(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n364_));
  INV_X1    g0172(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g0173(.A1(G69gat), .A2(G324gat), .ZN(new_n366_));
  AOI22_X1  g0174(.A1(new_n265_), .A2(new_n314_), .B1(new_n316_), .B2(new_n323_), .ZN(new_n367_));
  INV_X1    g0175(.A(new_n367_), .ZN(new_n368_));
  AND2_X1   g0176(.A1(G120gat), .A2(G273gat), .ZN(new_n369_));
  NOR2_X1   g0177(.A1(new_n309_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g0178(.A1(G103gat), .A2(G120gat), .A3(G273gat), .A4(G290gat), .ZN(new_n371_));
  INV_X1    g0179(.A(new_n371_), .ZN(new_n372_));
  OAI21_X1  g0180(.A(new_n310_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g0181(.A1(new_n309_), .A2(new_n371_), .A3(G86gat), .A4(G273gat), .ZN(new_n374_));
  NAND2_X1  g0182(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g0183(.A1(G86gat), .A2(G307gat), .ZN(new_n376_));
  INV_X1    g0184(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n378_));
  NOR2_X1   g0186(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g0187(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g0188(.A1(new_n368_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g0189(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g0190(.A(new_n376_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n383_));
  AND2_X1   g0191(.A1(G103gat), .A2(G273gat), .ZN(new_n384_));
  AND2_X1   g0192(.A1(G120gat), .A2(G290gat), .ZN(new_n385_));
  NAND2_X1  g0193(.A1(G120gat), .A2(G273gat), .ZN(new_n386_));
  AOI22_X1  g0194(.A1(new_n384_), .A2(new_n385_), .B1(new_n308_), .B2(new_n386_), .ZN(new_n387_));
  NOR3_X1   g0195(.A1(new_n308_), .A2(new_n312_), .A3(new_n194_), .ZN(new_n388_));
  OAI211_X1 g0196(.A(new_n374_), .B(new_n376_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  INV_X1    g0197(.A(new_n389_), .ZN(new_n390_));
  OAI21_X1  g0198(.A(new_n378_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g0199(.A1(new_n382_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g0200(.A(new_n367_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n393_));
  AOI21_X1  g0201(.A(new_n366_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g0202(.A1(new_n375_), .A2(new_n377_), .ZN(new_n395_));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n395_), .B2(new_n389_), .ZN(new_n396_));
  OAI211_X1 g0204(.A(new_n366_), .B(new_n393_), .C1(new_n396_), .C2(new_n381_), .ZN(new_n397_));
  INV_X1    g0205(.A(new_n397_), .ZN(new_n398_));
  OAI21_X1  g0206(.A(new_n365_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g0207(.A1(new_n214_), .A2(new_n261_), .ZN(new_n400_));
  INV_X1    g0208(.A(new_n400_), .ZN(new_n401_));
  OAI21_X1  g0209(.A(new_n393_), .B1(new_n396_), .B2(new_n381_), .ZN(new_n402_));
  NAND3_X1  g0210(.A1(new_n402_), .A2(G69gat), .A3(G324gat), .ZN(new_n403_));
  NAND3_X1  g0211(.A1(new_n403_), .A2(new_n364_), .A3(new_n397_), .ZN(new_n404_));
  NAND3_X1  g0212(.A1(new_n399_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g0213(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g0214(.A(new_n401_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g0215(.A(new_n363_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g0216(.A(new_n408_), .ZN(new_n409_));
  NOR3_X1   g0217(.A1(new_n363_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n410_));
  OAI21_X1  g0218(.A(new_n362_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g0219(.A(new_n363_), .ZN(new_n412_));
  INV_X1    g0220(.A(new_n407_), .ZN(new_n413_));
  NAND3_X1  g0221(.A1(new_n412_), .A2(new_n405_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g0222(.A(new_n362_), .ZN(new_n415_));
  NAND3_X1  g0223(.A1(new_n414_), .A2(new_n415_), .A3(new_n408_), .ZN(new_n416_));
  NAND2_X1  g0224(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g0225(.A1(new_n351_), .A2(new_n361_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g0226(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g0227(.A(new_n417_), .B1(new_n351_), .B2(new_n361_), .ZN(new_n420_));
  OAI21_X1  g0228(.A(new_n359_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g0229(.A(new_n420_), .ZN(new_n422_));
  INV_X1    g0230(.A(new_n359_), .ZN(new_n423_));
  NAND3_X1  g0231(.A1(new_n422_), .A2(new_n423_), .A3(new_n418_), .ZN(new_n424_));
  NAND2_X1  g0232(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g0233(.A(new_n354_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n426_));
  INV_X1    g0234(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g0235(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g0236(.A1(new_n426_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n429_));
  AND2_X1   g0237(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g0238(.A1(G1gat), .A2(G392gat), .ZN(new_n431_));
  XOR2_X1   g0239(.A(new_n431_), .B(KEYINPUT8), .Z(new_n432_));
  XNOR2_X1  g0240(.A(new_n430_), .B(new_n432_), .ZN(G3552gat));
  OR2_X1    g0241(.A1(new_n429_), .A2(KEYINPUT9), .ZN(new_n434_));
  NAND2_X1  g0242(.A1(new_n429_), .A2(KEYINPUT9), .ZN(new_n435_));
  NAND2_X1  g0243(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g0244(.A1(new_n428_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g0245(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g0246(.A(new_n422_), .B1(new_n419_), .B2(new_n359_), .ZN(new_n439_));
  NAND2_X1  g0247(.A1(new_n348_), .A2(G52gat), .ZN(new_n440_));
  INV_X1    g0248(.A(KEYINPUT11), .ZN(new_n441_));
  NAND2_X1  g0249(.A1(new_n405_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g0250(.A1(new_n312_), .A2(new_n232_), .ZN(new_n443_));
  INV_X1    g0251(.A(KEYINPUT12), .ZN(new_n444_));
  OAI21_X1  g0252(.A(new_n444_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n445_));
  OAI211_X1 g0253(.A(new_n310_), .B(KEYINPUT12), .C1(new_n370_), .C2(new_n372_), .ZN(new_n446_));
  AND3_X1   g0254(.A1(new_n389_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g0255(.A1(G120gat), .A2(G290gat), .ZN(new_n448_));
  NAND2_X1  g0256(.A1(G137gat), .A2(G273gat), .ZN(new_n449_));
  NAND2_X1  g0257(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g0258(.A1(G120gat), .A2(G137gat), .A3(G273gat), .A4(G290gat), .ZN(new_n451_));
  AOI22_X1  g0259(.A1(new_n450_), .A2(new_n451_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n452_));
  AND4_X1   g0260(.A1(G120gat), .A2(G137gat), .A3(G273gat), .A4(G290gat), .ZN(new_n453_));
  NOR2_X1   g0261(.A1(new_n453_), .A2(new_n371_), .ZN(new_n454_));
  INV_X1    g0262(.A(G103gat), .ZN(new_n455_));
  NOR2_X1   g0263(.A1(new_n455_), .A2(new_n245_), .ZN(new_n456_));
  NOR3_X1   g0264(.A1(new_n452_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g0265(.A(new_n456_), .ZN(new_n458_));
  AOI22_X1  g0266(.A1(G120gat), .A2(G290gat), .B1(G137gat), .B2(G273gat), .ZN(new_n459_));
  OAI21_X1  g0267(.A(new_n371_), .B1(new_n453_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g0268(.A1(new_n372_), .A2(new_n451_), .ZN(new_n461_));
  AOI21_X1  g0269(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g0270(.A(KEYINPUT13), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g0271(.A(new_n456_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n464_));
  NAND3_X1  g0272(.A1(new_n460_), .A2(new_n458_), .A3(new_n461_), .ZN(new_n465_));
  INV_X1    g0273(.A(KEYINPUT13), .ZN(new_n466_));
  NAND3_X1  g0274(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g0275(.A(new_n447_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g0276(.A(new_n466_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n469_));
  NAND3_X1  g0277(.A1(new_n389_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n470_));
  NOR2_X1   g0278(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g0279(.A(new_n443_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g0280(.A(KEYINPUT14), .ZN(new_n473_));
  AND3_X1   g0281(.A1(new_n464_), .A2(new_n466_), .A3(new_n465_), .ZN(new_n474_));
  OAI21_X1  g0282(.A(new_n470_), .B1(new_n474_), .B2(new_n469_), .ZN(new_n475_));
  NAND2_X1  g0283(.A1(new_n463_), .A2(new_n447_), .ZN(new_n476_));
  INV_X1    g0284(.A(new_n443_), .ZN(new_n477_));
  NAND3_X1  g0285(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND3_X1  g0286(.A1(new_n472_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n479_));
  NAND4_X1  g0287(.A1(new_n475_), .A2(KEYINPUT14), .A3(new_n477_), .A4(new_n476_), .ZN(new_n480_));
  NAND2_X1  g0288(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI22_X1  g0289(.A1(new_n382_), .A2(new_n391_), .B1(new_n366_), .B2(new_n393_), .ZN(new_n482_));
  NAND2_X1  g0290(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g0291(.A1(new_n318_), .A2(new_n261_), .ZN(new_n484_));
  INV_X1    g0292(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g0293(.A(new_n482_), .B1(new_n472_), .B2(new_n478_), .ZN(new_n486_));
  INV_X1    g0294(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g0295(.A1(new_n483_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g0296(.A(new_n482_), .ZN(new_n489_));
  AOI21_X1  g0297(.A(new_n489_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n490_));
  OAI21_X1  g0298(.A(new_n484_), .B1(new_n490_), .B2(new_n486_), .ZN(new_n491_));
  NAND3_X1  g0299(.A1(new_n442_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g0300(.A(KEYINPUT10), .ZN(new_n493_));
  NAND2_X1  g0301(.A1(new_n404_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g0302(.A1(new_n403_), .A2(new_n364_), .A3(KEYINPUT10), .A4(new_n397_), .ZN(new_n495_));
  AND2_X1   g0303(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g0304(.A1(new_n492_), .A2(new_n405_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g0305(.A1(new_n496_), .A2(new_n405_), .ZN(new_n498_));
  NAND4_X1  g0306(.A1(new_n498_), .A2(new_n442_), .A3(new_n488_), .A4(new_n491_), .ZN(new_n499_));
  AOI21_X1  g0307(.A(new_n440_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g0308(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g0309(.A(new_n410_), .B1(new_n415_), .B2(new_n408_), .ZN(new_n502_));
  INV_X1    g0310(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g0311(.A1(new_n497_), .A2(new_n499_), .A3(new_n440_), .ZN(new_n504_));
  NAND3_X1  g0312(.A1(new_n501_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g0313(.A(new_n504_), .ZN(new_n506_));
  OAI21_X1  g0314(.A(new_n502_), .B1(new_n506_), .B2(new_n500_), .ZN(new_n507_));
  NOR2_X1   g0315(.A1(new_n213_), .A2(new_n356_), .ZN(new_n508_));
  INV_X1    g0316(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g0317(.A1(new_n505_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g0318(.A(new_n503_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n511_));
  NOR3_X1   g0319(.A1(new_n506_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n512_));
  OAI21_X1  g0320(.A(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g0321(.A1(new_n439_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g0322(.A1(new_n513_), .A2(new_n510_), .ZN(new_n515_));
  OAI211_X1 g0323(.A(new_n515_), .B(new_n422_), .C1(new_n359_), .C2(new_n419_), .ZN(new_n516_));
  NAND2_X1  g0324(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g0325(.A1(G18gat), .A2(G392gat), .ZN(new_n518_));
  XOR2_X1   g0326(.A(new_n518_), .B(KEYINPUT15), .Z(new_n519_));
  OR2_X1    g0327(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g0328(.A1(new_n517_), .A2(new_n519_), .ZN(new_n521_));
  NAND3_X1  g0329(.A1(new_n438_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g0330(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  NAND2_X1  g0331(.A1(new_n430_), .A2(new_n432_), .ZN(new_n524_));
  NAND3_X1  g0332(.A1(new_n523_), .A2(new_n524_), .A3(new_n436_), .ZN(new_n525_));
  NAND2_X1  g0333(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g0334(.A1(G1gat), .A2(G409gat), .ZN(new_n527_));
  XNOR2_X1  g0335(.A(new_n526_), .B(new_n527_), .ZN(G3895gat));
  AOI22_X1  g0336(.A1(new_n526_), .A2(new_n527_), .B1(new_n438_), .B2(new_n523_), .ZN(new_n529_));
  NAND2_X1  g0337(.A1(new_n517_), .A2(KEYINPUT16), .ZN(new_n530_));
  INV_X1    g0338(.A(KEYINPUT16), .ZN(new_n531_));
  NAND3_X1  g0339(.A1(new_n514_), .A2(new_n516_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g0340(.A1(new_n530_), .A2(new_n519_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g0341(.A(new_n512_), .B1(new_n509_), .B2(new_n507_), .ZN(new_n534_));
  NAND3_X1  g0342(.A1(new_n498_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n535_));
  NAND2_X1  g0343(.A1(new_n504_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g0344(.A1(new_n455_), .A2(new_n232_), .ZN(new_n537_));
  INV_X1    g0345(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g0346(.A(G120gat), .ZN(new_n539_));
  NOR2_X1   g0347(.A1(new_n539_), .A2(new_n245_), .ZN(new_n540_));
  NAND2_X1  g0348(.A1(G137gat), .A2(G290gat), .ZN(new_n541_));
  NAND2_X1  g0349(.A1(G154gat), .A2(G273gat), .ZN(new_n542_));
  NAND2_X1  g0350(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g0351(.A1(G137gat), .A2(G154gat), .A3(G273gat), .A4(G290gat), .ZN(new_n544_));
  AND2_X1   g0352(.A1(G137gat), .A2(G290gat), .ZN(new_n545_));
  AOI22_X1  g0353(.A1(new_n543_), .A2(new_n544_), .B1(new_n369_), .B2(new_n545_), .ZN(new_n546_));
  AND4_X1   g0354(.A1(G137gat), .A2(G154gat), .A3(G273gat), .A4(G290gat), .ZN(new_n547_));
  NOR2_X1   g0355(.A1(new_n547_), .A2(new_n451_), .ZN(new_n548_));
  OAI21_X1  g0356(.A(new_n540_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  AOI22_X1  g0357(.A1(G137gat), .A2(G290gat), .B1(G154gat), .B2(G273gat), .ZN(new_n550_));
  OAI21_X1  g0358(.A(new_n451_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g0359(.A(new_n540_), .ZN(new_n552_));
  NAND2_X1  g0360(.A1(new_n453_), .A2(new_n544_), .ZN(new_n553_));
  NAND3_X1  g0361(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g0362(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g0363(.A(new_n460_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n556_));
  NAND2_X1  g0364(.A1(new_n556_), .A2(KEYINPUT17), .ZN(new_n557_));
  INV_X1    g0365(.A(KEYINPUT17), .ZN(new_n558_));
  OAI211_X1 g0366(.A(new_n460_), .B(new_n558_), .C1(new_n456_), .C2(new_n454_), .ZN(new_n559_));
  AOI21_X1  g0367(.A(new_n555_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  AND2_X1   g0368(.A1(new_n555_), .A2(new_n559_), .ZN(new_n561_));
  OAI21_X1  g0369(.A(new_n538_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g0370(.A1(new_n557_), .A2(new_n559_), .ZN(new_n563_));
  INV_X1    g0371(.A(new_n555_), .ZN(new_n564_));
  NAND2_X1  g0372(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g0373(.A1(new_n555_), .A2(new_n559_), .ZN(new_n566_));
  NAND3_X1  g0374(.A1(new_n565_), .A2(new_n537_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g0375(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g0376(.A(new_n477_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n569_));
  NOR3_X1   g0377(.A1(new_n447_), .A2(new_n457_), .A3(new_n462_), .ZN(new_n570_));
  INV_X1    g0378(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g0379(.A1(new_n568_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g0380(.A(new_n443_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n573_));
  OAI211_X1 g0381(.A(new_n562_), .B(new_n567_), .C1(new_n573_), .C2(new_n570_), .ZN(new_n574_));
  NOR2_X1   g0382(.A1(new_n312_), .A2(new_n261_), .ZN(new_n575_));
  INV_X1    g0383(.A(new_n575_), .ZN(new_n576_));
  AND3_X1   g0384(.A1(new_n572_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g0385(.A(new_n576_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n578_));
  NOR2_X1   g0386(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR3_X1   g0387(.A1(new_n490_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n580_));
  NOR2_X1   g0388(.A1(new_n481_), .A2(new_n482_), .ZN(new_n581_));
  OAI21_X1  g0389(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g0390(.A1(new_n572_), .A2(new_n574_), .ZN(new_n583_));
  NAND2_X1  g0391(.A1(new_n583_), .A2(new_n575_), .ZN(new_n584_));
  NAND3_X1  g0392(.A1(new_n572_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n585_));
  NAND2_X1  g0393(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g0394(.A(new_n581_), .ZN(new_n587_));
  NAND3_X1  g0395(.A1(new_n586_), .A2(new_n488_), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g0396(.A1(new_n302_), .A2(new_n318_), .ZN(new_n589_));
  INV_X1    g0397(.A(new_n589_), .ZN(new_n590_));
  AND3_X1   g0398(.A1(new_n582_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g0399(.A(new_n590_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n592_));
  NOR2_X1   g0400(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g0401(.A1(new_n536_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g0402(.A1(new_n214_), .A2(new_n356_), .ZN(new_n595_));
  INV_X1    g0403(.A(new_n595_), .ZN(new_n596_));
  OAI211_X1 g0404(.A(new_n504_), .B(new_n535_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n597_));
  NAND3_X1  g0405(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g0406(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g0407(.A(new_n596_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n600_));
  OAI21_X1  g0408(.A(new_n534_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g0409(.A1(new_n594_), .A2(new_n597_), .ZN(new_n602_));
  NAND2_X1  g0410(.A1(new_n602_), .A2(new_n595_), .ZN(new_n603_));
  OAI21_X1  g0411(.A(new_n505_), .B1(new_n511_), .B2(new_n508_), .ZN(new_n604_));
  NAND3_X1  g0412(.A1(new_n603_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n605_));
  NAND2_X1  g0413(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g0414(.A1(G35gat), .A2(G392gat), .ZN(new_n607_));
  XOR2_X1   g0415(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g0416(.A(KEYINPUT18), .ZN(new_n609_));
  NAND2_X1  g0417(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g0418(.A1(new_n606_), .A2(KEYINPUT18), .A3(new_n607_), .ZN(new_n611_));
  NAND4_X1  g0419(.A1(new_n533_), .A2(new_n514_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n612_));
  NAND3_X1  g0420(.A1(new_n514_), .A2(G18gat), .A3(G392gat), .ZN(new_n613_));
  NAND3_X1  g0421(.A1(new_n608_), .A2(new_n516_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g0422(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g0423(.A(G409gat), .ZN(new_n616_));
  NOR3_X1   g0424(.A1(new_n615_), .A2(new_n196_), .A3(new_n616_), .ZN(new_n617_));
  AOI22_X1  g0425(.A1(new_n612_), .A2(new_n614_), .B1(G18gat), .B2(G409gat), .ZN(new_n618_));
  NOR3_X1   g0426(.A1(new_n529_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g0427(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g0428(.A(new_n529_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n621_));
  NAND2_X1  g0429(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g0430(.A1(G1gat), .A2(G426gat), .ZN(new_n623_));
  XNOR2_X1  g0431(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g0432(.A(new_n624_), .B(KEYINPUT19), .Z(G4241gat));
  AOI21_X1  g0433(.A(new_n619_), .B1(new_n623_), .B2(new_n621_), .ZN(new_n626_));
  OAI21_X1  g0434(.A(new_n615_), .B1(new_n196_), .B2(new_n616_), .ZN(new_n627_));
  NAND2_X1  g0435(.A1(new_n610_), .A2(new_n611_), .ZN(new_n628_));
  NAND2_X1  g0436(.A1(new_n613_), .A2(new_n516_), .ZN(new_n629_));
  NOR2_X1   g0437(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g0438(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g0439(.A1(new_n601_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n632_));
  INV_X1    g0440(.A(KEYINPUT29), .ZN(new_n633_));
  NAND2_X1  g0441(.A1(new_n603_), .A2(new_n598_), .ZN(new_n634_));
  INV_X1    g0442(.A(KEYINPUT20), .ZN(new_n635_));
  AOI21_X1  g0443(.A(new_n534_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g0444(.A1(new_n603_), .A2(KEYINPUT20), .A3(new_n598_), .ZN(new_n637_));
  AOI22_X1  g0445(.A1(new_n632_), .A2(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g0446(.A1(new_n601_), .A2(new_n605_), .A3(KEYINPUT29), .A4(new_n607_), .ZN(new_n639_));
  NAND2_X1  g0447(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g0448(.A1(G69gat), .A2(G375gat), .ZN(new_n641_));
  XOR2_X1   g0449(.A(new_n641_), .B(KEYINPUT28), .Z(new_n642_));
  INV_X1    g0450(.A(new_n642_), .ZN(new_n643_));
  INV_X1    g0451(.A(new_n574_), .ZN(new_n644_));
  AOI21_X1  g0452(.A(new_n644_), .B1(new_n576_), .B2(new_n572_), .ZN(new_n645_));
  NAND2_X1  g0453(.A1(new_n565_), .A2(new_n566_), .ZN(new_n646_));
  AOI22_X1  g0454(.A1(new_n646_), .A2(new_n538_), .B1(new_n564_), .B2(new_n556_), .ZN(new_n647_));
  INV_X1    g0455(.A(G137gat), .ZN(new_n648_));
  NOR2_X1   g0456(.A1(new_n648_), .A2(new_n245_), .ZN(new_n649_));
  INV_X1    g0457(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g0458(.A1(G154gat), .A2(G290gat), .ZN(new_n651_));
  NAND2_X1  g0459(.A1(G171gat), .A2(G273gat), .ZN(new_n652_));
  NAND2_X1  g0460(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g0461(.A1(G154gat), .A2(G171gat), .A3(G273gat), .A4(G290gat), .ZN(new_n654_));
  AND2_X1   g0462(.A1(G137gat), .A2(G273gat), .ZN(new_n655_));
  AND2_X1   g0463(.A1(G154gat), .A2(G290gat), .ZN(new_n656_));
  AOI22_X1  g0464(.A1(new_n653_), .A2(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AND4_X1   g0465(.A1(G154gat), .A2(G171gat), .A3(G273gat), .A4(G290gat), .ZN(new_n658_));
  NOR2_X1   g0466(.A1(new_n658_), .A2(new_n544_), .ZN(new_n659_));
  OAI21_X1  g0467(.A(new_n650_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  AOI22_X1  g0468(.A1(G154gat), .A2(G290gat), .B1(G171gat), .B2(G273gat), .ZN(new_n661_));
  OAI21_X1  g0469(.A(new_n544_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g0470(.A1(new_n547_), .A2(new_n654_), .ZN(new_n663_));
  NAND3_X1  g0471(.A1(new_n662_), .A2(new_n649_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g0472(.A1(new_n660_), .A2(new_n664_), .A3(KEYINPUT25), .ZN(new_n665_));
  NOR3_X1   g0473(.A1(new_n657_), .A2(new_n659_), .A3(new_n650_), .ZN(new_n666_));
  INV_X1    g0474(.A(KEYINPUT25), .ZN(new_n667_));
  NAND2_X1  g0475(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g0476(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g0477(.A(new_n546_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n670_));
  INV_X1    g0478(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g0479(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g0480(.A1(new_n539_), .A2(new_n232_), .ZN(new_n673_));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n674_));
  NAND2_X1  g0482(.A1(new_n551_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g0483(.A1(new_n546_), .A2(KEYINPUT26), .ZN(new_n676_));
  AND2_X1   g0484(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g0485(.A(new_n649_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n678_));
  OAI211_X1 g0486(.A(new_n677_), .B(new_n554_), .C1(new_n666_), .C2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g0487(.A1(new_n672_), .A2(new_n673_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g0488(.A(new_n673_), .ZN(new_n681_));
  AOI21_X1  g0489(.A(new_n670_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n682_));
  NOR2_X1   g0490(.A1(new_n666_), .A2(new_n678_), .ZN(new_n683_));
  NAND3_X1  g0491(.A1(new_n554_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n684_));
  NOR2_X1   g0492(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g0493(.A(new_n681_), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g0494(.A1(new_n680_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g0495(.A(KEYINPUT24), .B1(new_n646_), .B2(new_n538_), .ZN(new_n688_));
  OAI21_X1  g0496(.A(new_n647_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g0497(.A1(new_n564_), .A2(new_n556_), .ZN(new_n690_));
  NAND2_X1  g0498(.A1(new_n562_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g0499(.A(KEYINPUT24), .ZN(new_n692_));
  NAND2_X1  g0500(.A1(new_n562_), .A2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g0501(.A1(new_n691_), .A2(new_n693_), .A3(new_n686_), .A4(new_n680_), .ZN(new_n694_));
  NOR2_X1   g0502(.A1(new_n455_), .A2(new_n261_), .ZN(new_n695_));
  INV_X1    g0503(.A(new_n695_), .ZN(new_n696_));
  AND3_X1   g0504(.A1(new_n689_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g0505(.A(new_n696_), .B1(new_n689_), .B2(new_n694_), .ZN(new_n698_));
  OAI21_X1  g0506(.A(new_n645_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g0507(.A1(new_n689_), .A2(new_n694_), .ZN(new_n700_));
  NAND2_X1  g0508(.A1(new_n700_), .A2(new_n695_), .ZN(new_n701_));
  NAND2_X1  g0509(.A1(new_n585_), .A2(new_n574_), .ZN(new_n702_));
  NAND3_X1  g0510(.A1(new_n689_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n703_));
  NAND3_X1  g0511(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NOR2_X1   g0512(.A1(new_n302_), .A2(new_n312_), .ZN(new_n705_));
  INV_X1    g0513(.A(new_n705_), .ZN(new_n706_));
  AND3_X1   g0514(.A1(new_n699_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g0515(.A(new_n706_), .B1(new_n699_), .B2(new_n704_), .ZN(new_n708_));
  NOR2_X1   g0516(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g0517(.A1(new_n699_), .A2(new_n704_), .ZN(new_n710_));
  NAND2_X1  g0518(.A1(new_n710_), .A2(new_n706_), .ZN(new_n711_));
  NAND2_X1  g0519(.A1(new_n711_), .A2(KEYINPUT27), .ZN(new_n712_));
  NAND3_X1  g0520(.A1(new_n582_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n713_));
  OAI21_X1  g0521(.A(KEYINPUT23), .B1(new_n580_), .B2(new_n581_), .ZN(new_n714_));
  INV_X1    g0522(.A(KEYINPUT23), .ZN(new_n715_));
  NAND3_X1  g0523(.A1(new_n488_), .A2(new_n715_), .A3(new_n587_), .ZN(new_n716_));
  NAND3_X1  g0524(.A1(new_n714_), .A2(new_n716_), .A3(new_n579_), .ZN(new_n717_));
  NAND2_X1  g0525(.A1(new_n713_), .A2(new_n717_), .ZN(new_n718_));
  AND3_X1   g0526(.A1(new_n709_), .A2(new_n712_), .A3(new_n718_), .ZN(new_n719_));
  NAND3_X1  g0527(.A1(new_n699_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n720_));
  INV_X1    g0528(.A(new_n708_), .ZN(new_n721_));
  AOI22_X1  g0529(.A1(new_n712_), .A2(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g0530(.A(new_n643_), .B1(new_n719_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g0531(.A1(new_n721_), .A2(new_n720_), .ZN(new_n724_));
  AND2_X1   g0532(.A1(new_n713_), .A2(new_n717_), .ZN(new_n725_));
  INV_X1    g0533(.A(KEYINPUT27), .ZN(new_n726_));
  AOI21_X1  g0534(.A(new_n726_), .B1(new_n710_), .B2(new_n706_), .ZN(new_n727_));
  OAI21_X1  g0535(.A(new_n724_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g0536(.A1(new_n709_), .A2(new_n712_), .A3(new_n718_), .ZN(new_n729_));
  NAND3_X1  g0537(.A1(new_n728_), .A2(new_n642_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g0538(.A1(new_n594_), .A2(KEYINPUT22), .ZN(new_n731_));
  NAND3_X1  g0539(.A1(new_n723_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g0540(.A(new_n597_), .ZN(new_n733_));
  OAI21_X1  g0541(.A(new_n594_), .B1(new_n733_), .B2(new_n595_), .ZN(new_n734_));
  INV_X1    g0542(.A(new_n734_), .ZN(new_n735_));
  NAND2_X1  g0543(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g0544(.A1(new_n734_), .A2(new_n723_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n737_));
  NAND2_X1  g0545(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g0546(.A1(new_n738_), .A2(G52gat), .A3(G392gat), .ZN(new_n739_));
  NAND2_X1  g0547(.A1(G52gat), .A2(G392gat), .ZN(new_n740_));
  NAND3_X1  g0548(.A1(new_n736_), .A2(new_n740_), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g0549(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g0550(.A1(new_n640_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g0551(.A(new_n635_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n744_));
  NAND3_X1  g0552(.A1(new_n744_), .A2(new_n637_), .A3(new_n604_), .ZN(new_n745_));
  NAND2_X1  g0553(.A1(new_n745_), .A2(KEYINPUT21), .ZN(new_n746_));
  INV_X1    g0554(.A(KEYINPUT21), .ZN(new_n747_));
  NAND4_X1  g0555(.A1(new_n744_), .A2(new_n637_), .A3(new_n747_), .A4(new_n604_), .ZN(new_n748_));
  NAND3_X1  g0556(.A1(new_n746_), .A2(new_n632_), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g0557(.A(new_n743_), .B1(new_n742_), .B2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g0558(.A1(new_n213_), .A2(new_n616_), .ZN(new_n751_));
  INV_X1    g0559(.A(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g0560(.A(new_n750_), .B(new_n752_), .ZN(new_n753_));
  NAND3_X1  g0561(.A1(new_n627_), .A2(new_n631_), .A3(new_n753_), .ZN(new_n754_));
  NAND2_X1  g0562(.A1(G18gat), .A2(G426gat), .ZN(new_n755_));
  XNOR2_X1  g0563(.A(new_n750_), .B(new_n751_), .ZN(new_n756_));
  OAI21_X1  g0564(.A(new_n756_), .B1(new_n618_), .B2(new_n630_), .ZN(new_n757_));
  NAND3_X1  g0565(.A1(new_n754_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g0566(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g0567(.A(new_n755_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n760_));
  OAI21_X1  g0568(.A(new_n626_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g0569(.A(new_n761_), .ZN(new_n762_));
  NOR3_X1   g0570(.A1(new_n626_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n763_));
  NOR2_X1   g0571(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g0572(.A(G443gat), .ZN(new_n765_));
  NOR2_X1   g0573(.A1(new_n193_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g0574(.A(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g0575(.A(new_n764_), .B(new_n767_), .ZN(G4591gat));
  OR2_X1    g0576(.A1(new_n756_), .A2(KEYINPUT30), .ZN(new_n769_));
  NAND2_X1  g0577(.A1(new_n627_), .A2(new_n631_), .ZN(new_n770_));
  NAND2_X1  g0578(.A1(new_n756_), .A2(KEYINPUT30), .ZN(new_n771_));
  NAND3_X1  g0579(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g0580(.A1(new_n758_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g0581(.A(G426gat), .ZN(new_n774_));
  NOR2_X1   g0582(.A1(new_n213_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g0583(.A(new_n775_), .ZN(new_n776_));
  NOR2_X1   g0584(.A1(new_n742_), .A2(new_n749_), .ZN(new_n777_));
  AOI22_X1  g0585(.A1(new_n638_), .A2(new_n639_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n778_));
  OAI21_X1  g0586(.A(new_n752_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g0587(.A(KEYINPUT37), .ZN(new_n780_));
  NAND2_X1  g0588(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g0589(.A(KEYINPUT37), .B(new_n752_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g0590(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g0591(.A(new_n742_), .B1(new_n639_), .B2(new_n638_), .ZN(new_n784_));
  INV_X1    g0592(.A(new_n784_), .ZN(new_n785_));
  NOR2_X1   g0593(.A1(new_n214_), .A2(new_n616_), .ZN(new_n786_));
  INV_X1    g0594(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g0595(.A1(new_n734_), .A2(new_n723_), .A3(new_n730_), .ZN(new_n788_));
  NAND2_X1  g0596(.A1(new_n741_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g0597(.A1(new_n709_), .A2(new_n718_), .ZN(new_n790_));
  NAND2_X1  g0598(.A1(new_n730_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g0599(.A1(new_n312_), .A2(new_n356_), .ZN(new_n792_));
  NAND3_X1  g0600(.A1(new_n691_), .A2(new_n686_), .A3(new_n680_), .ZN(new_n793_));
  NAND2_X1  g0601(.A1(new_n703_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g0602(.A(KEYINPUT33), .ZN(new_n795_));
  NOR2_X1   g0603(.A1(new_n648_), .A2(new_n232_), .ZN(new_n796_));
  NAND3_X1  g0604(.A1(KEYINPUT32), .A2(G154gat), .A3(G307gat), .ZN(new_n797_));
  NAND2_X1  g0605(.A1(G171gat), .A2(G290gat), .ZN(new_n798_));
  NAND2_X1  g0606(.A1(G188gat), .A2(G273gat), .ZN(new_n799_));
  NAND2_X1  g0607(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g0608(.A1(G171gat), .A2(G188gat), .A3(G273gat), .A4(G290gat), .ZN(new_n801_));
  INV_X1    g0609(.A(new_n542_), .ZN(new_n802_));
  AND2_X1   g0610(.A1(G171gat), .A2(G290gat), .ZN(new_n803_));
  AOI22_X1  g0611(.A1(new_n800_), .A2(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AND4_X1   g0612(.A1(G171gat), .A2(G188gat), .A3(G273gat), .A4(G290gat), .ZN(new_n805_));
  NOR2_X1   g0613(.A1(new_n805_), .A2(new_n654_), .ZN(new_n806_));
  OAI21_X1  g0614(.A(new_n797_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g0615(.A(new_n663_), .B1(new_n657_), .B2(new_n650_), .ZN(new_n808_));
  AOI22_X1  g0616(.A1(G171gat), .A2(G290gat), .B1(G188gat), .B2(G273gat), .ZN(new_n809_));
  OAI21_X1  g0617(.A(new_n654_), .B1(new_n805_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g0618(.A1(new_n658_), .A2(new_n801_), .ZN(new_n811_));
  NAND2_X1  g0619(.A1(G154gat), .A2(G307gat), .ZN(new_n812_));
  INV_X1    g0620(.A(KEYINPUT32), .ZN(new_n813_));
  NAND2_X1  g0621(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g0622(.A1(new_n814_), .A2(new_n797_), .ZN(new_n815_));
  NAND3_X1  g0623(.A1(new_n810_), .A2(new_n811_), .A3(new_n815_), .ZN(new_n816_));
  AND3_X1   g0624(.A1(new_n807_), .A2(new_n808_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g0625(.A(new_n808_), .B1(new_n816_), .B2(new_n807_), .ZN(new_n818_));
  OAI21_X1  g0626(.A(new_n796_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g0627(.A(new_n659_), .B1(new_n662_), .B2(new_n649_), .ZN(new_n820_));
  AND3_X1   g0628(.A1(new_n810_), .A2(new_n811_), .A3(new_n815_), .ZN(new_n821_));
  INV_X1    g0629(.A(new_n797_), .ZN(new_n822_));
  AOI21_X1  g0630(.A(new_n822_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n823_));
  OAI21_X1  g0631(.A(new_n820_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g0632(.A(new_n796_), .ZN(new_n825_));
  NAND3_X1  g0633(.A1(new_n807_), .A2(new_n808_), .A3(new_n816_), .ZN(new_n826_));
  NAND3_X1  g0634(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g0635(.A1(new_n819_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g0636(.A1(new_n665_), .A2(new_n668_), .A3(new_n684_), .ZN(new_n829_));
  AND3_X1   g0637(.A1(new_n828_), .A2(new_n686_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g0638(.A(new_n828_), .B1(new_n686_), .B2(new_n829_), .ZN(new_n831_));
  OAI21_X1  g0639(.A(new_n795_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g0640(.A1(new_n539_), .A2(new_n261_), .ZN(new_n833_));
  NAND2_X1  g0641(.A1(new_n686_), .A2(new_n829_), .ZN(new_n834_));
  AND2_X1   g0642(.A1(new_n819_), .A2(new_n827_), .ZN(new_n835_));
  NAND2_X1  g0643(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g0644(.A1(new_n828_), .A2(new_n686_), .A3(new_n829_), .ZN(new_n837_));
  NAND3_X1  g0645(.A1(new_n836_), .A2(KEYINPUT33), .A3(new_n837_), .ZN(new_n838_));
  NAND3_X1  g0646(.A1(new_n832_), .A2(new_n833_), .A3(new_n838_), .ZN(new_n839_));
  NOR3_X1   g0647(.A1(new_n830_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n840_));
  INV_X1    g0648(.A(new_n840_), .ZN(new_n841_));
  NAND3_X1  g0649(.A1(new_n794_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g0650(.A1(new_n348_), .A2(G103gat), .ZN(new_n843_));
  INV_X1    g0651(.A(new_n833_), .ZN(new_n844_));
  AOI21_X1  g0652(.A(new_n844_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n845_));
  OAI211_X1 g0653(.A(new_n703_), .B(new_n793_), .C1(new_n840_), .C2(new_n845_), .ZN(new_n846_));
  AND3_X1   g0654(.A1(new_n842_), .A2(new_n843_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g0655(.A(new_n843_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n848_));
  OAI21_X1  g0656(.A(KEYINPUT34), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g0657(.A(KEYINPUT31), .ZN(new_n850_));
  NAND2_X1  g0658(.A1(new_n704_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g0659(.A1(new_n701_), .A2(new_n702_), .A3(KEYINPUT31), .A4(new_n703_), .ZN(new_n852_));
  NAND3_X1  g0660(.A1(new_n720_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g0661(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g0662(.A1(new_n842_), .A2(new_n846_), .ZN(new_n855_));
  INV_X1    g0663(.A(KEYINPUT34), .ZN(new_n856_));
  NAND3_X1  g0664(.A1(new_n855_), .A2(new_n856_), .A3(new_n843_), .ZN(new_n857_));
  NAND3_X1  g0665(.A1(new_n849_), .A2(new_n854_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g0666(.A(new_n853_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n859_));
  AOI21_X1  g0667(.A(new_n792_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g0668(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g0669(.A1(new_n858_), .A2(new_n792_), .A3(new_n859_), .ZN(new_n862_));
  NAND3_X1  g0670(.A1(new_n791_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AND3_X1   g0671(.A1(new_n858_), .A2(new_n792_), .A3(new_n859_), .ZN(new_n864_));
  OAI211_X1 g0672(.A(new_n730_), .B(new_n790_), .C1(new_n864_), .C2(new_n860_), .ZN(new_n865_));
  NAND2_X1  g0673(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g0674(.A(G392gat), .ZN(new_n867_));
  NOR2_X1   g0675(.A1(new_n318_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g0676(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g0677(.A(new_n868_), .ZN(new_n870_));
  NAND3_X1  g0678(.A1(new_n863_), .A2(new_n865_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g0679(.A(KEYINPUT35), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g0680(.A1(new_n863_), .A2(new_n865_), .A3(KEYINPUT35), .ZN(new_n873_));
  INV_X1    g0681(.A(new_n873_), .ZN(new_n874_));
  OAI211_X1 g0682(.A(KEYINPUT36), .B(new_n789_), .C1(new_n872_), .C2(new_n874_), .ZN(new_n875_));
  AND3_X1   g0683(.A1(new_n863_), .A2(new_n865_), .A3(new_n870_), .ZN(new_n876_));
  AOI21_X1  g0684(.A(new_n870_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n877_));
  NOR3_X1   g0685(.A1(new_n789_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g0686(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g0687(.A1(new_n875_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g0688(.A(KEYINPUT35), .ZN(new_n881_));
  OAI21_X1  g0689(.A(new_n881_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n882_));
  NAND2_X1  g0690(.A1(new_n882_), .A2(new_n873_), .ZN(new_n883_));
  AOI21_X1  g0691(.A(KEYINPUT36), .B1(new_n883_), .B2(new_n789_), .ZN(new_n884_));
  OAI21_X1  g0692(.A(new_n787_), .B1(new_n880_), .B2(new_n884_), .ZN(new_n885_));
  AND2_X1   g0693(.A1(new_n741_), .A2(new_n788_), .ZN(new_n886_));
  AOI21_X1  g0694(.A(new_n886_), .B1(new_n882_), .B2(new_n873_), .ZN(new_n887_));
  AOI21_X1  g0695(.A(new_n878_), .B1(new_n887_), .B2(KEYINPUT36), .ZN(new_n888_));
  OAI21_X1  g0696(.A(new_n789_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n889_));
  INV_X1    g0697(.A(KEYINPUT36), .ZN(new_n890_));
  NAND2_X1  g0698(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g0699(.A1(new_n888_), .A2(new_n786_), .A3(new_n891_), .ZN(new_n892_));
  AOI22_X1  g0700(.A1(new_n783_), .A2(new_n785_), .B1(new_n885_), .B2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g0701(.A(new_n784_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n894_));
  AND3_X1   g0702(.A1(new_n894_), .A2(new_n885_), .A3(new_n892_), .ZN(new_n895_));
  OAI21_X1  g0703(.A(new_n776_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g0704(.A1(new_n894_), .A2(new_n885_), .A3(new_n892_), .ZN(new_n897_));
  NOR3_X1   g0705(.A1(new_n880_), .A2(new_n884_), .A3(new_n787_), .ZN(new_n898_));
  AOI21_X1  g0706(.A(new_n786_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n899_));
  NOR2_X1   g0707(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g0708(.A(new_n784_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n901_));
  OAI21_X1  g0709(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  OR2_X1    g0710(.A1(new_n902_), .A2(new_n776_), .ZN(new_n903_));
  NAND3_X1  g0711(.A1(new_n773_), .A2(new_n896_), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g0712(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g0713(.A(new_n773_), .B1(new_n896_), .B2(new_n903_), .ZN(new_n906_));
  NOR2_X1   g0714(.A1(new_n196_), .A2(new_n765_), .ZN(new_n907_));
  AND2_X1   g0715(.A1(new_n907_), .A2(KEYINPUT38), .ZN(new_n908_));
  NOR2_X1   g0716(.A1(new_n907_), .A2(KEYINPUT38), .ZN(new_n909_));
  OAI22_X1  g0717(.A1(new_n905_), .A2(new_n906_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g0718(.A1(new_n903_), .A2(new_n896_), .ZN(new_n911_));
  NAND3_X1  g0719(.A1(new_n911_), .A2(new_n758_), .A3(new_n772_), .ZN(new_n912_));
  OAI211_X1 g0720(.A(new_n912_), .B(new_n904_), .C1(KEYINPUT38), .C2(new_n907_), .ZN(new_n913_));
  AND2_X1   g0721(.A1(new_n910_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1  g0722(.A(new_n763_), .B1(new_n767_), .B2(new_n761_), .ZN(new_n915_));
  XOR2_X1   g0723(.A(new_n914_), .B(new_n915_), .Z(new_n916_));
  NAND2_X1  g0724(.A1(G1gat), .A2(G460gat), .ZN(new_n917_));
  XNOR2_X1  g0725(.A(new_n916_), .B(new_n917_), .ZN(G4946gat));
  AOI21_X1  g0726(.A(new_n915_), .B1(new_n910_), .B2(new_n913_), .ZN(new_n919_));
  NAND2_X1  g0727(.A1(new_n914_), .A2(new_n915_), .ZN(new_n920_));
  AOI21_X1  g0728(.A(new_n919_), .B1(new_n920_), .B2(new_n917_), .ZN(new_n921_));
  NOR2_X1   g0729(.A1(new_n213_), .A2(new_n765_), .ZN(new_n922_));
  NAND2_X1  g0730(.A1(new_n885_), .A2(new_n892_), .ZN(new_n923_));
  NOR2_X1   g0731(.A1(new_n901_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g0732(.A(new_n924_), .ZN(new_n925_));
  NAND2_X1  g0733(.A1(new_n896_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g0734(.A1(new_n873_), .A2(new_n870_), .ZN(new_n927_));
  AOI21_X1  g0735(.A(KEYINPUT35), .B1(new_n863_), .B2(new_n865_), .ZN(new_n928_));
  OAI21_X1  g0736(.A(KEYINPUT39), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g0737(.A1(new_n866_), .A2(new_n881_), .ZN(new_n930_));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n931_));
  NAND4_X1  g0739(.A1(new_n930_), .A2(new_n931_), .A3(new_n873_), .A4(new_n870_), .ZN(new_n932_));
  NOR2_X1   g0740(.A1(new_n312_), .A2(new_n867_), .ZN(new_n933_));
  NAND3_X1  g0741(.A1(new_n842_), .A2(new_n843_), .A3(new_n846_), .ZN(new_n934_));
  NOR2_X1   g0742(.A1(new_n840_), .A2(new_n845_), .ZN(new_n935_));
  NAND2_X1  g0743(.A1(new_n935_), .A2(new_n794_), .ZN(new_n936_));
  NAND2_X1  g0744(.A1(new_n934_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g0745(.A1(new_n648_), .A2(new_n261_), .ZN(new_n938_));
  NAND2_X1  g0746(.A1(new_n827_), .A2(new_n824_), .ZN(new_n939_));
  OAI21_X1  g0747(.A(new_n811_), .B1(new_n804_), .B2(new_n812_), .ZN(new_n940_));
  NAND2_X1  g0748(.A1(G188gat), .A2(G290gat), .ZN(new_n941_));
  INV_X1    g0749(.A(G205gat), .ZN(new_n942_));
  OAI21_X1  g0750(.A(new_n941_), .B1(new_n942_), .B2(new_n194_), .ZN(new_n943_));
  NAND4_X1  g0751(.A1(G188gat), .A2(G205gat), .A3(G273gat), .A4(G290gat), .ZN(new_n944_));
  AOI21_X1  g0752(.A(new_n805_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  INV_X1    g0753(.A(G171gat), .ZN(new_n946_));
  NOR2_X1   g0754(.A1(new_n946_), .A2(new_n245_), .ZN(new_n947_));
  AND4_X1   g0755(.A1(G188gat), .A2(G205gat), .A3(G273gat), .A4(G290gat), .ZN(new_n948_));
  NOR2_X1   g0756(.A1(new_n948_), .A2(new_n801_), .ZN(new_n949_));
  NOR3_X1   g0757(.A1(new_n945_), .A2(new_n947_), .A3(new_n949_), .ZN(new_n950_));
  INV_X1    g0758(.A(new_n947_), .ZN(new_n951_));
  AOI22_X1  g0759(.A1(G188gat), .A2(G290gat), .B1(G205gat), .B2(G273gat), .ZN(new_n952_));
  OAI21_X1  g0760(.A(new_n801_), .B1(new_n948_), .B2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g0761(.A1(new_n805_), .A2(new_n944_), .ZN(new_n954_));
  AOI21_X1  g0762(.A(new_n951_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  OAI21_X1  g0763(.A(new_n940_), .B1(new_n950_), .B2(new_n955_), .ZN(new_n956_));
  INV_X1    g0764(.A(G154gat), .ZN(new_n957_));
  NOR2_X1   g0765(.A1(new_n957_), .A2(new_n232_), .ZN(new_n958_));
  INV_X1    g0766(.A(new_n958_), .ZN(new_n959_));
  OAI21_X1  g0767(.A(new_n947_), .B1(new_n945_), .B2(new_n949_), .ZN(new_n960_));
  INV_X1    g0768(.A(new_n812_), .ZN(new_n961_));
  AOI21_X1  g0769(.A(new_n806_), .B1(new_n810_), .B2(new_n961_), .ZN(new_n962_));
  NAND3_X1  g0770(.A1(new_n953_), .A2(new_n951_), .A3(new_n954_), .ZN(new_n963_));
  NAND3_X1  g0771(.A1(new_n960_), .A2(new_n962_), .A3(new_n963_), .ZN(new_n964_));
  NAND3_X1  g0772(.A1(new_n956_), .A2(new_n959_), .A3(new_n964_), .ZN(new_n965_));
  AOI21_X1  g0773(.A(new_n959_), .B1(new_n956_), .B2(new_n964_), .ZN(new_n966_));
  INV_X1    g0774(.A(new_n966_), .ZN(new_n967_));
  AOI21_X1  g0775(.A(new_n939_), .B1(new_n965_), .B2(new_n967_), .ZN(new_n968_));
  INV_X1    g0776(.A(new_n965_), .ZN(new_n969_));
  AOI21_X1  g0777(.A(new_n818_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n970_));
  NOR3_X1   g0778(.A1(new_n969_), .A2(new_n970_), .A3(new_n966_), .ZN(new_n971_));
  OAI21_X1  g0779(.A(new_n938_), .B1(new_n968_), .B2(new_n971_), .ZN(new_n972_));
  NAND3_X1  g0780(.A1(new_n967_), .A2(new_n939_), .A3(new_n965_), .ZN(new_n973_));
  OAI21_X1  g0781(.A(new_n970_), .B1(new_n969_), .B2(new_n966_), .ZN(new_n974_));
  INV_X1    g0782(.A(new_n938_), .ZN(new_n975_));
  NAND3_X1  g0783(.A1(new_n973_), .A2(new_n974_), .A3(new_n975_), .ZN(new_n976_));
  NAND2_X1  g0784(.A1(new_n972_), .A2(new_n976_), .ZN(new_n977_));
  OAI21_X1  g0785(.A(new_n836_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n978_));
  NAND2_X1  g0786(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  AOI21_X1  g0787(.A(new_n833_), .B1(new_n832_), .B2(new_n838_), .ZN(new_n980_));
  NAND3_X1  g0788(.A1(new_n972_), .A2(new_n976_), .A3(new_n836_), .ZN(new_n981_));
  OAI21_X1  g0789(.A(new_n979_), .B1(new_n980_), .B2(new_n981_), .ZN(new_n982_));
  NOR2_X1   g0790(.A1(new_n302_), .A2(new_n539_), .ZN(new_n983_));
  INV_X1    g0791(.A(new_n983_), .ZN(new_n984_));
  NAND2_X1  g0792(.A1(new_n982_), .A2(new_n984_), .ZN(new_n985_));
  OAI211_X1 g0793(.A(new_n979_), .B(new_n983_), .C1(new_n980_), .C2(new_n981_), .ZN(new_n986_));
  NAND3_X1  g0794(.A1(new_n937_), .A2(new_n985_), .A3(new_n986_), .ZN(new_n987_));
  AND3_X1   g0795(.A1(new_n836_), .A2(KEYINPUT33), .A3(new_n837_), .ZN(new_n988_));
  AOI21_X1  g0796(.A(KEYINPUT33), .B1(new_n836_), .B2(new_n837_), .ZN(new_n989_));
  OAI21_X1  g0797(.A(new_n844_), .B1(new_n988_), .B2(new_n989_), .ZN(new_n990_));
  INV_X1    g0798(.A(new_n981_), .ZN(new_n991_));
  NAND2_X1  g0799(.A1(new_n990_), .A2(new_n991_), .ZN(new_n992_));
  AOI21_X1  g0800(.A(new_n983_), .B1(new_n992_), .B2(new_n979_), .ZN(new_n993_));
  INV_X1    g0801(.A(new_n986_), .ZN(new_n994_));
  OAI211_X1 g0802(.A(new_n934_), .B(new_n936_), .C1(new_n993_), .C2(new_n994_), .ZN(new_n995_));
  NAND2_X1  g0803(.A1(new_n987_), .A2(new_n995_), .ZN(new_n996_));
  NOR2_X1   g0804(.A1(new_n455_), .A2(new_n356_), .ZN(new_n997_));
  NAND2_X1  g0805(.A1(new_n996_), .A2(new_n997_), .ZN(new_n998_));
  INV_X1    g0806(.A(new_n997_), .ZN(new_n999_));
  NAND3_X1  g0807(.A1(new_n987_), .A2(new_n995_), .A3(new_n999_), .ZN(new_n1000_));
  NAND2_X1  g0808(.A1(new_n998_), .A2(new_n1000_), .ZN(new_n1001_));
  INV_X1    g0809(.A(KEYINPUT40), .ZN(new_n1002_));
  NAND2_X1  g0810(.A1(new_n853_), .A2(new_n1002_), .ZN(new_n1003_));
  NAND4_X1  g0811(.A1(new_n720_), .A2(KEYINPUT40), .A3(new_n851_), .A4(new_n852_), .ZN(new_n1004_));
  NAND4_X1  g0812(.A1(new_n1003_), .A2(new_n849_), .A3(new_n857_), .A4(new_n1004_), .ZN(new_n1005_));
  AOI21_X1  g0813(.A(new_n1001_), .B1(new_n861_), .B2(new_n1005_), .ZN(new_n1006_));
  AND3_X1   g0814(.A1(new_n987_), .A2(new_n995_), .A3(new_n999_), .ZN(new_n1007_));
  AOI21_X1  g0815(.A(new_n999_), .B1(new_n987_), .B2(new_n995_), .ZN(new_n1008_));
  NOR2_X1   g0816(.A1(new_n1007_), .A2(new_n1008_), .ZN(new_n1009_));
  INV_X1    g0817(.A(new_n1005_), .ZN(new_n1010_));
  NOR3_X1   g0818(.A1(new_n1009_), .A2(new_n860_), .A3(new_n1010_), .ZN(new_n1011_));
  OAI21_X1  g0819(.A(new_n933_), .B1(new_n1006_), .B2(new_n1011_), .ZN(new_n1012_));
  NAND3_X1  g0820(.A1(new_n861_), .A2(new_n1001_), .A3(new_n1005_), .ZN(new_n1013_));
  OAI21_X1  g0821(.A(new_n1009_), .B1(new_n860_), .B2(new_n1010_), .ZN(new_n1014_));
  INV_X1    g0822(.A(new_n933_), .ZN(new_n1015_));
  NAND3_X1  g0823(.A1(new_n1013_), .A2(new_n1014_), .A3(new_n1015_), .ZN(new_n1016_));
  AND3_X1   g0824(.A1(new_n1012_), .A2(new_n863_), .A3(new_n1016_), .ZN(new_n1017_));
  NAND3_X1  g0825(.A1(new_n929_), .A2(new_n932_), .A3(new_n1017_), .ZN(new_n1018_));
  NOR2_X1   g0826(.A1(new_n318_), .A2(new_n616_), .ZN(new_n1019_));
  NAND2_X1  g0827(.A1(new_n1012_), .A2(new_n1016_), .ZN(new_n1020_));
  NAND2_X1  g0828(.A1(new_n871_), .A2(new_n863_), .ZN(new_n1021_));
  NAND2_X1  g0829(.A1(new_n1020_), .A2(new_n1021_), .ZN(new_n1022_));
  AND3_X1   g0830(.A1(new_n1018_), .A2(new_n1019_), .A3(new_n1022_), .ZN(new_n1023_));
  AOI21_X1  g0831(.A(new_n1019_), .B1(new_n1018_), .B2(new_n1022_), .ZN(new_n1024_));
  NOR2_X1   g0832(.A1(new_n1023_), .A2(new_n1024_), .ZN(new_n1025_));
  NOR3_X1   g0833(.A1(new_n886_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n1026_));
  OAI21_X1  g0834(.A(new_n1025_), .B1(new_n899_), .B2(new_n1026_), .ZN(new_n1027_));
  NAND2_X1  g0835(.A1(new_n1018_), .A2(new_n1022_), .ZN(new_n1028_));
  INV_X1    g0836(.A(new_n1019_), .ZN(new_n1029_));
  NAND2_X1  g0837(.A1(new_n1028_), .A2(new_n1029_), .ZN(new_n1030_));
  NAND3_X1  g0838(.A1(new_n1018_), .A2(new_n1019_), .A3(new_n1022_), .ZN(new_n1031_));
  NAND2_X1  g0839(.A1(new_n1030_), .A2(new_n1031_), .ZN(new_n1032_));
  INV_X1    g0840(.A(new_n1026_), .ZN(new_n1033_));
  NAND3_X1  g0841(.A1(new_n1032_), .A2(new_n885_), .A3(new_n1033_), .ZN(new_n1034_));
  NOR2_X1   g0842(.A1(new_n214_), .A2(new_n774_), .ZN(new_n1035_));
  INV_X1    g0843(.A(new_n1035_), .ZN(new_n1036_));
  AND3_X1   g0844(.A1(new_n1027_), .A2(new_n1034_), .A3(new_n1036_), .ZN(new_n1037_));
  AOI21_X1  g0845(.A(new_n1036_), .B1(new_n1027_), .B2(new_n1034_), .ZN(new_n1038_));
  NOR2_X1   g0846(.A1(new_n1037_), .A2(new_n1038_), .ZN(new_n1039_));
  NOR2_X1   g0847(.A1(new_n926_), .A2(new_n1039_), .ZN(new_n1040_));
  NAND2_X1  g0848(.A1(new_n1027_), .A2(new_n1034_), .ZN(new_n1041_));
  NAND2_X1  g0849(.A1(new_n1041_), .A2(new_n1035_), .ZN(new_n1042_));
  NAND3_X1  g0850(.A1(new_n1027_), .A2(new_n1034_), .A3(new_n1036_), .ZN(new_n1043_));
  NAND2_X1  g0851(.A1(new_n1042_), .A2(new_n1043_), .ZN(new_n1044_));
  AOI21_X1  g0852(.A(new_n924_), .B1(new_n902_), .B2(new_n776_), .ZN(new_n1045_));
  NOR2_X1   g0853(.A1(new_n1044_), .A2(new_n1045_), .ZN(new_n1046_));
  OAI21_X1  g0854(.A(new_n922_), .B1(new_n1040_), .B2(new_n1046_), .ZN(new_n1047_));
  NAND2_X1  g0855(.A1(new_n926_), .A2(new_n1039_), .ZN(new_n1048_));
  NAND2_X1  g0856(.A1(new_n1044_), .A2(new_n1045_), .ZN(new_n1049_));
  INV_X1    g0857(.A(new_n922_), .ZN(new_n1050_));
  NAND3_X1  g0858(.A1(new_n1048_), .A2(new_n1049_), .A3(new_n1050_), .ZN(new_n1051_));
  AND2_X1   g0859(.A1(new_n1047_), .A2(new_n1051_), .ZN(new_n1052_));
  OAI21_X1  g0860(.A(new_n904_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n1053_));
  OR2_X1    g0861(.A1(new_n1052_), .A2(new_n1053_), .ZN(new_n1054_));
  INV_X1    g0862(.A(G460gat), .ZN(new_n1055_));
  NOR2_X1   g0863(.A1(new_n196_), .A2(new_n1055_), .ZN(new_n1056_));
  NAND3_X1  g0864(.A1(new_n1053_), .A2(new_n1051_), .A3(new_n1047_), .ZN(new_n1057_));
  AND3_X1   g0865(.A1(new_n1054_), .A2(new_n1056_), .A3(new_n1057_), .ZN(new_n1058_));
  AOI21_X1  g0866(.A(new_n1056_), .B1(new_n1054_), .B2(new_n1057_), .ZN(new_n1059_));
  OAI21_X1  g0867(.A(new_n921_), .B1(new_n1058_), .B2(new_n1059_), .ZN(new_n1060_));
  INV_X1    g0868(.A(KEYINPUT41), .ZN(new_n1061_));
  NAND2_X1  g0869(.A1(new_n1060_), .A2(new_n1061_), .ZN(new_n1062_));
  OAI211_X1 g0870(.A(new_n921_), .B(KEYINPUT41), .C1(new_n1058_), .C2(new_n1059_), .ZN(new_n1063_));
  NAND3_X1  g0871(.A1(new_n1054_), .A2(new_n1056_), .A3(new_n1057_), .ZN(new_n1064_));
  XNOR2_X1  g0872(.A(new_n1064_), .B(KEYINPUT42), .ZN(new_n1065_));
  NOR2_X1   g0873(.A1(new_n921_), .A2(new_n1059_), .ZN(new_n1066_));
  AOI22_X1  g0874(.A1(new_n1062_), .A2(new_n1063_), .B1(new_n1065_), .B2(new_n1066_), .ZN(new_n1067_));
  NAND2_X1  g0875(.A1(G1gat), .A2(G477gat), .ZN(new_n1068_));
  XOR2_X1   g0876(.A(new_n1068_), .B(KEYINPUT43), .Z(new_n1069_));
  INV_X1    g0877(.A(new_n1069_), .ZN(new_n1070_));
  XNOR2_X1  g0878(.A(new_n1067_), .B(new_n1070_), .ZN(G5308gat));
  NAND2_X1  g0879(.A1(new_n1057_), .A2(new_n1056_), .ZN(new_n1072_));
  AND2_X1   g0880(.A1(new_n1054_), .A2(new_n1072_), .ZN(new_n1073_));
  AOI21_X1  g0881(.A(new_n1046_), .B1(new_n1050_), .B2(new_n1049_), .ZN(new_n1074_));
  AOI21_X1  g0882(.A(new_n971_), .B1(new_n975_), .B2(new_n974_), .ZN(new_n1075_));
  AOI21_X1  g0883(.A(new_n962_), .B1(new_n960_), .B2(new_n963_), .ZN(new_n1076_));
  OAI21_X1  g0884(.A(new_n964_), .B1(new_n1076_), .B2(new_n958_), .ZN(new_n1077_));
  INV_X1    g0885(.A(KEYINPUT46), .ZN(new_n1078_));
  NAND2_X1  g0886(.A1(new_n1077_), .A2(new_n1078_), .ZN(new_n1079_));
  OAI211_X1 g0887(.A(KEYINPUT46), .B(new_n964_), .C1(new_n1076_), .C2(new_n958_), .ZN(new_n1080_));
  NAND2_X1  g0888(.A1(new_n1079_), .A2(new_n1080_), .ZN(new_n1081_));
  AOI21_X1  g0889(.A(new_n945_), .B1(new_n951_), .B2(new_n954_), .ZN(new_n1082_));
  NAND2_X1  g0890(.A1(G205gat), .A2(G290gat), .ZN(new_n1083_));
  NAND2_X1  g0891(.A1(G222gat), .A2(G273gat), .ZN(new_n1084_));
  NAND2_X1  g0892(.A1(new_n1083_), .A2(new_n1084_), .ZN(new_n1085_));
  NAND4_X1  g0893(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1086_));
  INV_X1    g0894(.A(new_n799_), .ZN(new_n1087_));
  AND2_X1   g0895(.A1(G205gat), .A2(G290gat), .ZN(new_n1088_));
  AOI22_X1  g0896(.A1(new_n1085_), .A2(new_n1086_), .B1(new_n1087_), .B2(new_n1088_), .ZN(new_n1089_));
  AND4_X1   g0897(.A1(G205gat), .A2(G222gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1090_));
  NOR2_X1   g0898(.A1(new_n1090_), .A2(new_n944_), .ZN(new_n1091_));
  INV_X1    g0899(.A(G188gat), .ZN(new_n1092_));
  NOR2_X1   g0900(.A1(new_n1092_), .A2(new_n245_), .ZN(new_n1093_));
  INV_X1    g0901(.A(new_n1093_), .ZN(new_n1094_));
  NOR3_X1   g0902(.A1(new_n1089_), .A2(new_n1091_), .A3(new_n1094_), .ZN(new_n1095_));
  INV_X1    g0903(.A(KEYINPUT45), .ZN(new_n1096_));
  OAI21_X1  g0904(.A(new_n1094_), .B1(new_n1089_), .B2(new_n1091_), .ZN(new_n1097_));
  AOI21_X1  g0905(.A(new_n1095_), .B1(new_n1096_), .B2(new_n1097_), .ZN(new_n1098_));
  OAI211_X1 g0906(.A(KEYINPUT45), .B(new_n1094_), .C1(new_n1089_), .C2(new_n1091_), .ZN(new_n1099_));
  AOI21_X1  g0907(.A(new_n1082_), .B1(new_n1098_), .B2(new_n1099_), .ZN(new_n1100_));
  NOR2_X1   g0908(.A1(new_n946_), .A2(new_n232_), .ZN(new_n1101_));
  NAND2_X1  g0909(.A1(new_n1085_), .A2(new_n1086_), .ZN(new_n1102_));
  NAND2_X1  g0910(.A1(new_n1102_), .A2(new_n944_), .ZN(new_n1103_));
  NAND2_X1  g0911(.A1(new_n948_), .A2(new_n1086_), .ZN(new_n1104_));
  NAND3_X1  g0912(.A1(new_n1103_), .A2(new_n1093_), .A3(new_n1104_), .ZN(new_n1105_));
  AND3_X1   g0913(.A1(new_n1082_), .A2(new_n1097_), .A3(new_n1105_), .ZN(new_n1106_));
  NOR3_X1   g0914(.A1(new_n1100_), .A2(new_n1101_), .A3(new_n1106_), .ZN(new_n1107_));
  INV_X1    g0915(.A(new_n1101_), .ZN(new_n1108_));
  NAND2_X1  g0916(.A1(new_n1097_), .A2(new_n1096_), .ZN(new_n1109_));
  NAND3_X1  g0917(.A1(new_n1109_), .A2(new_n1099_), .A3(new_n1105_), .ZN(new_n1110_));
  INV_X1    g0918(.A(new_n1082_), .ZN(new_n1111_));
  NAND2_X1  g0919(.A1(new_n1110_), .A2(new_n1111_), .ZN(new_n1112_));
  INV_X1    g0920(.A(new_n1106_), .ZN(new_n1113_));
  AOI21_X1  g0921(.A(new_n1108_), .B1(new_n1112_), .B2(new_n1113_), .ZN(new_n1114_));
  OAI21_X1  g0922(.A(new_n1081_), .B1(new_n1107_), .B2(new_n1114_), .ZN(new_n1115_));
  NOR2_X1   g0923(.A1(new_n957_), .A2(new_n261_), .ZN(new_n1116_));
  OAI21_X1  g0924(.A(new_n1101_), .B1(new_n1100_), .B2(new_n1106_), .ZN(new_n1117_));
  NAND3_X1  g0925(.A1(new_n1112_), .A2(new_n1113_), .A3(new_n1108_), .ZN(new_n1118_));
  NAND3_X1  g0926(.A1(new_n1117_), .A2(new_n1118_), .A3(new_n1079_), .ZN(new_n1119_));
  AND3_X1   g0927(.A1(new_n1115_), .A2(new_n1116_), .A3(new_n1119_), .ZN(new_n1120_));
  AOI21_X1  g0928(.A(new_n1116_), .B1(new_n1115_), .B2(new_n1119_), .ZN(new_n1121_));
  OAI21_X1  g0929(.A(new_n1075_), .B1(new_n1120_), .B2(new_n1121_), .ZN(new_n1122_));
  AND3_X1   g0930(.A1(new_n1117_), .A2(new_n1118_), .A3(new_n1079_), .ZN(new_n1123_));
  AOI22_X1  g0931(.A1(new_n1117_), .A2(new_n1118_), .B1(new_n1080_), .B2(new_n1079_), .ZN(new_n1124_));
  OAI22_X1  g0932(.A1(new_n1123_), .A2(new_n1124_), .B1(new_n957_), .B2(new_n261_), .ZN(new_n1125_));
  INV_X1    g0933(.A(new_n1075_), .ZN(new_n1126_));
  NAND3_X1  g0934(.A1(new_n1115_), .A2(new_n1116_), .A3(new_n1119_), .ZN(new_n1127_));
  NAND3_X1  g0935(.A1(new_n1125_), .A2(new_n1126_), .A3(new_n1127_), .ZN(new_n1128_));
  OAI211_X1 g0936(.A(new_n1122_), .B(new_n1128_), .C1(new_n648_), .C2(new_n302_), .ZN(new_n1129_));
  NOR2_X1   g0937(.A1(new_n302_), .A2(new_n648_), .ZN(new_n1130_));
  NOR3_X1   g0938(.A1(new_n1120_), .A2(new_n1121_), .A3(new_n1075_), .ZN(new_n1131_));
  AOI21_X1  g0939(.A(new_n1126_), .B1(new_n1125_), .B2(new_n1127_), .ZN(new_n1132_));
  OAI21_X1  g0940(.A(new_n1130_), .B1(new_n1131_), .B2(new_n1132_), .ZN(new_n1133_));
  AOI21_X1  g0941(.A(new_n977_), .B1(new_n841_), .B2(new_n836_), .ZN(new_n1134_));
  OAI211_X1 g0942(.A(new_n1129_), .B(new_n1133_), .C1(new_n993_), .C2(new_n1134_), .ZN(new_n1135_));
  NAND2_X1  g0943(.A1(new_n1133_), .A2(new_n1129_), .ZN(new_n1136_));
  AOI21_X1  g0944(.A(new_n1134_), .B1(new_n982_), .B2(new_n984_), .ZN(new_n1137_));
  NAND2_X1  g0945(.A1(new_n1136_), .A2(new_n1137_), .ZN(new_n1138_));
  NOR2_X1   g0946(.A1(new_n539_), .A2(new_n356_), .ZN(new_n1139_));
  XOR2_X1   g0947(.A(new_n1139_), .B(KEYINPUT47), .Z(new_n1140_));
  AND3_X1   g0948(.A1(new_n1135_), .A2(new_n1138_), .A3(new_n1140_), .ZN(new_n1141_));
  AOI21_X1  g0949(.A(new_n1140_), .B1(new_n1135_), .B2(new_n1138_), .ZN(new_n1142_));
  OAI211_X1 g0950(.A(new_n987_), .B(new_n1000_), .C1(new_n1141_), .C2(new_n1142_), .ZN(new_n1143_));
  AOI21_X1  g0951(.A(new_n937_), .B1(new_n985_), .B2(new_n986_), .ZN(new_n1144_));
  OAI21_X1  g0952(.A(new_n987_), .B1(new_n1144_), .B2(new_n997_), .ZN(new_n1145_));
  NAND2_X1  g0953(.A1(new_n1135_), .A2(new_n1138_), .ZN(new_n1146_));
  INV_X1    g0954(.A(new_n1140_), .ZN(new_n1147_));
  NAND2_X1  g0955(.A1(new_n1146_), .A2(new_n1147_), .ZN(new_n1148_));
  OAI211_X1 g0956(.A(new_n1135_), .B(new_n1138_), .C1(new_n539_), .C2(new_n356_), .ZN(new_n1149_));
  NAND3_X1  g0957(.A1(new_n1145_), .A2(new_n1148_), .A3(new_n1149_), .ZN(new_n1150_));
  NOR2_X1   g0958(.A1(new_n455_), .A2(new_n867_), .ZN(new_n1151_));
  INV_X1    g0959(.A(new_n1151_), .ZN(new_n1152_));
  AND3_X1   g0960(.A1(new_n1143_), .A2(new_n1150_), .A3(new_n1152_), .ZN(new_n1153_));
  AOI21_X1  g0961(.A(new_n1152_), .B1(new_n1143_), .B2(new_n1150_), .ZN(new_n1154_));
  OAI211_X1 g0962(.A(new_n1016_), .B(new_n1014_), .C1(new_n1153_), .C2(new_n1154_), .ZN(new_n1155_));
  NOR2_X1   g0963(.A1(new_n1153_), .A2(new_n1154_), .ZN(new_n1156_));
  OAI21_X1  g0964(.A(new_n1014_), .B1(new_n1011_), .B2(new_n933_), .ZN(new_n1157_));
  NAND2_X1  g0965(.A1(new_n1156_), .A2(new_n1157_), .ZN(new_n1158_));
  NOR2_X1   g0966(.A1(new_n312_), .A2(new_n616_), .ZN(new_n1159_));
  INV_X1    g0967(.A(new_n1159_), .ZN(new_n1160_));
  AND3_X1   g0968(.A1(new_n1155_), .A2(new_n1158_), .A3(new_n1160_), .ZN(new_n1161_));
  AOI21_X1  g0969(.A(new_n1160_), .B1(new_n1155_), .B2(new_n1158_), .ZN(new_n1162_));
  OAI21_X1  g0970(.A(KEYINPUT48), .B1(new_n1161_), .B2(new_n1162_), .ZN(new_n1163_));
  AOI21_X1  g0971(.A(new_n1020_), .B1(new_n863_), .B2(new_n871_), .ZN(new_n1164_));
  INV_X1    g0972(.A(new_n1164_), .ZN(new_n1165_));
  NAND2_X1  g0973(.A1(new_n1155_), .A2(new_n1158_), .ZN(new_n1166_));
  INV_X1    g0974(.A(KEYINPUT48), .ZN(new_n1167_));
  NAND3_X1  g0975(.A1(new_n1166_), .A2(new_n1167_), .A3(new_n1160_), .ZN(new_n1168_));
  AND3_X1   g0976(.A1(new_n1163_), .A2(new_n1165_), .A3(new_n1168_), .ZN(new_n1169_));
  INV_X1    g0977(.A(KEYINPUT44), .ZN(new_n1170_));
  INV_X1    g0978(.A(new_n1022_), .ZN(new_n1171_));
  NAND3_X1  g0979(.A1(new_n1012_), .A2(new_n863_), .A3(new_n1016_), .ZN(new_n1172_));
  NAND3_X1  g0980(.A1(new_n930_), .A2(new_n873_), .A3(new_n870_), .ZN(new_n1173_));
  AOI21_X1  g0981(.A(new_n1172_), .B1(new_n1173_), .B2(KEYINPUT39), .ZN(new_n1174_));
  AOI21_X1  g0982(.A(new_n1171_), .B1(new_n1174_), .B2(new_n932_), .ZN(new_n1175_));
  OAI21_X1  g0983(.A(new_n1170_), .B1(new_n1175_), .B2(new_n1019_), .ZN(new_n1176_));
  NAND2_X1  g0984(.A1(new_n1024_), .A2(KEYINPUT44), .ZN(new_n1177_));
  NAND3_X1  g0985(.A1(new_n1169_), .A2(new_n1176_), .A3(new_n1177_), .ZN(new_n1178_));
  OR2_X1    g0986(.A1(new_n1161_), .A2(new_n1162_), .ZN(new_n1179_));
  OAI21_X1  g0987(.A(new_n1179_), .B1(new_n1024_), .B2(new_n1164_), .ZN(new_n1180_));
  INV_X1    g0988(.A(KEYINPUT49), .ZN(new_n1181_));
  NAND2_X1  g0989(.A1(new_n1180_), .A2(new_n1181_), .ZN(new_n1182_));
  OAI211_X1 g0990(.A(KEYINPUT49), .B(new_n1179_), .C1(new_n1024_), .C2(new_n1164_), .ZN(new_n1183_));
  NAND3_X1  g0991(.A1(new_n1178_), .A2(new_n1182_), .A3(new_n1183_), .ZN(new_n1184_));
  NOR2_X1   g0992(.A1(new_n318_), .A2(new_n774_), .ZN(new_n1185_));
  INV_X1    g0993(.A(new_n1185_), .ZN(new_n1186_));
  NAND2_X1  g0994(.A1(new_n1184_), .A2(new_n1186_), .ZN(new_n1187_));
  NOR3_X1   g0995(.A1(new_n1025_), .A2(new_n899_), .A3(new_n1026_), .ZN(new_n1188_));
  OAI21_X1  g0996(.A(new_n1027_), .B1(new_n1188_), .B2(new_n1035_), .ZN(new_n1189_));
  NAND4_X1  g0997(.A1(new_n1178_), .A2(new_n1182_), .A3(new_n1185_), .A4(new_n1183_), .ZN(new_n1190_));
  AND3_X1   g0998(.A1(new_n1187_), .A2(new_n1189_), .A3(new_n1190_), .ZN(new_n1191_));
  AOI21_X1  g0999(.A(new_n1189_), .B1(new_n1187_), .B2(new_n1190_), .ZN(new_n1192_));
  NOR2_X1   g1000(.A1(new_n214_), .A2(new_n765_), .ZN(new_n1193_));
  NOR3_X1   g1001(.A1(new_n1191_), .A2(new_n1192_), .A3(new_n1193_), .ZN(new_n1194_));
  INV_X1    g1002(.A(new_n1193_), .ZN(new_n1195_));
  NAND2_X1  g1003(.A1(new_n1187_), .A2(new_n1190_), .ZN(new_n1196_));
  INV_X1    g1004(.A(new_n1189_), .ZN(new_n1197_));
  NAND2_X1  g1005(.A1(new_n1196_), .A2(new_n1197_), .ZN(new_n1198_));
  NAND3_X1  g1006(.A1(new_n1187_), .A2(new_n1189_), .A3(new_n1190_), .ZN(new_n1199_));
  AOI21_X1  g1007(.A(new_n1195_), .B1(new_n1198_), .B2(new_n1199_), .ZN(new_n1200_));
  OAI21_X1  g1008(.A(new_n1074_), .B1(new_n1194_), .B2(new_n1200_), .ZN(new_n1201_));
  OAI21_X1  g1009(.A(new_n1048_), .B1(new_n1040_), .B2(new_n922_), .ZN(new_n1202_));
  NAND3_X1  g1010(.A1(new_n1198_), .A2(new_n1195_), .A3(new_n1199_), .ZN(new_n1203_));
  OAI21_X1  g1011(.A(new_n1193_), .B1(new_n1191_), .B2(new_n1192_), .ZN(new_n1204_));
  NAND3_X1  g1012(.A1(new_n1202_), .A2(new_n1203_), .A3(new_n1204_), .ZN(new_n1205_));
  NOR2_X1   g1013(.A1(new_n213_), .A2(new_n1055_), .ZN(new_n1206_));
  INV_X1    g1014(.A(new_n1206_), .ZN(new_n1207_));
  NAND3_X1  g1015(.A1(new_n1201_), .A2(new_n1205_), .A3(new_n1207_), .ZN(new_n1208_));
  INV_X1    g1016(.A(new_n1208_), .ZN(new_n1209_));
  AOI21_X1  g1017(.A(new_n1207_), .B1(new_n1201_), .B2(new_n1205_), .ZN(new_n1210_));
  NOR2_X1   g1018(.A1(new_n1209_), .A2(new_n1210_), .ZN(new_n1211_));
  NAND2_X1  g1019(.A1(new_n1073_), .A2(new_n1211_), .ZN(new_n1212_));
  NAND2_X1  g1020(.A1(new_n1054_), .A2(new_n1072_), .ZN(new_n1213_));
  OAI21_X1  g1021(.A(new_n1213_), .B1(new_n1209_), .B2(new_n1210_), .ZN(new_n1214_));
  INV_X1    g1022(.A(G477gat), .ZN(new_n1215_));
  OAI211_X1 g1023(.A(new_n1212_), .B(new_n1214_), .C1(new_n196_), .C2(new_n1215_), .ZN(new_n1216_));
  NAND2_X1  g1024(.A1(new_n1212_), .A2(new_n1214_), .ZN(new_n1217_));
  NAND3_X1  g1025(.A1(new_n1217_), .A2(G18gat), .A3(G477gat), .ZN(new_n1218_));
  NAND2_X1  g1026(.A1(new_n1062_), .A2(new_n1063_), .ZN(new_n1219_));
  NAND2_X1  g1027(.A1(new_n1065_), .A2(new_n1066_), .ZN(new_n1220_));
  AOI21_X1  g1028(.A(new_n1070_), .B1(new_n1219_), .B2(new_n1220_), .ZN(new_n1221_));
  NOR2_X1   g1029(.A1(new_n1058_), .A2(new_n1059_), .ZN(new_n1222_));
  NOR2_X1   g1030(.A1(new_n1222_), .A2(new_n921_), .ZN(new_n1223_));
  OAI211_X1 g1031(.A(new_n1216_), .B(new_n1218_), .C1(new_n1221_), .C2(new_n1223_), .ZN(new_n1224_));
  INV_X1    g1032(.A(new_n1223_), .ZN(new_n1225_));
  NAND2_X1  g1033(.A1(new_n1218_), .A2(new_n1216_), .ZN(new_n1226_));
  OAI211_X1 g1034(.A(new_n1225_), .B(new_n1226_), .C1(new_n1067_), .C2(new_n1070_), .ZN(new_n1227_));
  NAND2_X1  g1035(.A1(new_n1224_), .A2(new_n1227_), .ZN(new_n1228_));
  NAND2_X1  g1036(.A1(G1gat), .A2(G494gat), .ZN(new_n1229_));
  XOR2_X1   g1037(.A(new_n1229_), .B(KEYINPUT50), .Z(new_n1230_));
  XOR2_X1   g1038(.A(new_n1228_), .B(new_n1230_), .Z(G5672gat));
  NAND3_X1  g1039(.A1(new_n1224_), .A2(G1gat), .A3(G494gat), .ZN(new_n1232_));
  INV_X1    g1040(.A(KEYINPUT51), .ZN(new_n1233_));
  NAND2_X1  g1041(.A1(new_n1212_), .A2(new_n1233_), .ZN(new_n1234_));
  NAND3_X1  g1042(.A1(new_n1073_), .A2(KEYINPUT51), .A3(new_n1211_), .ZN(new_n1235_));
  NAND3_X1  g1043(.A1(new_n1216_), .A2(new_n1234_), .A3(new_n1235_), .ZN(new_n1236_));
  INV_X1    g1044(.A(KEYINPUT52), .ZN(new_n1237_));
  OAI21_X1  g1045(.A(new_n1237_), .B1(new_n1194_), .B2(new_n1200_), .ZN(new_n1238_));
  NAND3_X1  g1046(.A1(new_n1204_), .A2(new_n1203_), .A3(KEYINPUT52), .ZN(new_n1239_));
  NAND3_X1  g1047(.A1(new_n1238_), .A2(new_n1202_), .A3(new_n1239_), .ZN(new_n1240_));
  NAND2_X1  g1048(.A1(new_n1208_), .A2(new_n1240_), .ZN(new_n1241_));
  OAI21_X1  g1049(.A(new_n1199_), .B1(new_n1192_), .B2(new_n1193_), .ZN(new_n1242_));
  INV_X1    g1050(.A(new_n1242_), .ZN(new_n1243_));
  NAND3_X1  g1051(.A1(new_n1143_), .A2(new_n1150_), .A3(new_n1152_), .ZN(new_n1244_));
  NAND3_X1  g1052(.A1(new_n1135_), .A2(new_n1138_), .A3(new_n1140_), .ZN(new_n1245_));
  NAND3_X1  g1053(.A1(new_n1145_), .A2(new_n1148_), .A3(new_n1245_), .ZN(new_n1246_));
  NAND2_X1  g1054(.A1(new_n1244_), .A2(new_n1246_), .ZN(new_n1247_));
  INV_X1    g1055(.A(new_n1247_), .ZN(new_n1248_));
  OAI21_X1  g1056(.A(KEYINPUT53), .B1(new_n993_), .B2(new_n1134_), .ZN(new_n1249_));
  INV_X1    g1057(.A(KEYINPUT53), .ZN(new_n1250_));
  NAND2_X1  g1058(.A1(new_n1137_), .A2(new_n1250_), .ZN(new_n1251_));
  NAND4_X1  g1059(.A1(new_n1249_), .A2(new_n1251_), .A3(new_n1129_), .A4(new_n1133_), .ZN(new_n1252_));
  NAND2_X1  g1060(.A1(new_n1149_), .A2(new_n1252_), .ZN(new_n1253_));
  INV_X1    g1061(.A(KEYINPUT54), .ZN(new_n1254_));
  NAND2_X1  g1062(.A1(new_n1125_), .A2(new_n1254_), .ZN(new_n1255_));
  NOR2_X1   g1063(.A1(new_n946_), .A2(new_n261_), .ZN(new_n1256_));
  NAND2_X1  g1064(.A1(new_n1118_), .A2(new_n1112_), .ZN(new_n1257_));
  INV_X1    g1065(.A(KEYINPUT56), .ZN(new_n1258_));
  NAND4_X1  g1066(.A1(G222gat), .A2(G239gat), .A3(G273gat), .A4(G290gat), .ZN(new_n1259_));
  NAND2_X1  g1067(.A1(new_n1090_), .A2(new_n1259_), .ZN(new_n1260_));
  AND2_X1   g1068(.A1(G222gat), .A2(G273gat), .ZN(new_n1261_));
  AND2_X1   g1069(.A1(G239gat), .A2(G290gat), .ZN(new_n1262_));
  NAND2_X1  g1070(.A1(G222gat), .A2(G290gat), .ZN(new_n1263_));
  NAND2_X1  g1071(.A1(G239gat), .A2(G273gat), .ZN(new_n1264_));
  AOI22_X1  g1072(.A1(new_n1261_), .A2(new_n1262_), .B1(new_n1263_), .B2(new_n1264_), .ZN(new_n1265_));
  OAI211_X1 g1073(.A(new_n1258_), .B(new_n1260_), .C1(new_n1265_), .C2(new_n1090_), .ZN(new_n1266_));
  NOR2_X1   g1074(.A1(new_n942_), .A2(new_n245_), .ZN(new_n1267_));
  INV_X1    g1075(.A(new_n1267_), .ZN(new_n1268_));
  NAND2_X1  g1076(.A1(new_n1263_), .A2(new_n1264_), .ZN(new_n1269_));
  NAND2_X1  g1077(.A1(new_n1269_), .A2(new_n1259_), .ZN(new_n1270_));
  OAI21_X1  g1078(.A(KEYINPUT56), .B1(new_n1270_), .B2(new_n1090_), .ZN(new_n1271_));
  NAND3_X1  g1079(.A1(new_n1266_), .A2(new_n1268_), .A3(new_n1271_), .ZN(new_n1272_));
  OAI211_X1 g1080(.A(new_n1267_), .B(new_n1260_), .C1(new_n1265_), .C2(new_n1090_), .ZN(new_n1273_));
  INV_X1    g1081(.A(KEYINPUT57), .ZN(new_n1274_));
  NAND2_X1  g1082(.A1(new_n1273_), .A2(new_n1274_), .ZN(new_n1275_));
  NAND2_X1  g1083(.A1(new_n1270_), .A2(new_n1086_), .ZN(new_n1276_));
  NAND4_X1  g1084(.A1(new_n1276_), .A2(KEYINPUT57), .A3(new_n1267_), .A4(new_n1260_), .ZN(new_n1277_));
  NAND3_X1  g1085(.A1(new_n1272_), .A2(new_n1275_), .A3(new_n1277_), .ZN(new_n1278_));
  AOI21_X1  g1086(.A(new_n1091_), .B1(new_n1103_), .B2(new_n1093_), .ZN(new_n1279_));
  NAND2_X1  g1087(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1280_));
  NOR2_X1   g1088(.A1(new_n1092_), .A2(new_n232_), .ZN(new_n1281_));
  INV_X1    g1089(.A(new_n1281_), .ZN(new_n1282_));
  NAND2_X1  g1090(.A1(new_n1266_), .A2(new_n1271_), .ZN(new_n1283_));
  NAND2_X1  g1091(.A1(new_n1283_), .A2(new_n1267_), .ZN(new_n1284_));
  INV_X1    g1092(.A(new_n1279_), .ZN(new_n1285_));
  NAND3_X1  g1093(.A1(new_n1284_), .A2(new_n1285_), .A3(new_n1272_), .ZN(new_n1286_));
  AND3_X1   g1094(.A1(new_n1280_), .A2(new_n1282_), .A3(new_n1286_), .ZN(new_n1287_));
  AOI21_X1  g1095(.A(new_n1282_), .B1(new_n1280_), .B2(new_n1286_), .ZN(new_n1288_));
  NOR2_X1   g1096(.A1(new_n1287_), .A2(new_n1288_), .ZN(new_n1289_));
  NAND2_X1  g1097(.A1(new_n1112_), .A2(KEYINPUT55), .ZN(new_n1290_));
  AOI21_X1  g1098(.A(new_n1257_), .B1(new_n1289_), .B2(new_n1290_), .ZN(new_n1291_));
  NAND2_X1  g1099(.A1(new_n1280_), .A2(new_n1286_), .ZN(new_n1292_));
  NAND2_X1  g1100(.A1(new_n1292_), .A2(new_n1281_), .ZN(new_n1293_));
  NAND3_X1  g1101(.A1(new_n1280_), .A2(new_n1282_), .A3(new_n1286_), .ZN(new_n1294_));
  AND4_X1   g1102(.A1(new_n1257_), .A2(new_n1293_), .A3(new_n1294_), .A4(new_n1290_), .ZN(new_n1295_));
  OAI21_X1  g1103(.A(new_n1256_), .B1(new_n1291_), .B2(new_n1295_), .ZN(new_n1296_));
  NAND3_X1  g1104(.A1(new_n1293_), .A2(new_n1294_), .A3(new_n1290_), .ZN(new_n1297_));
  INV_X1    g1105(.A(new_n1257_), .ZN(new_n1298_));
  NAND2_X1  g1106(.A1(new_n1297_), .A2(new_n1298_), .ZN(new_n1299_));
  INV_X1    g1107(.A(new_n1256_), .ZN(new_n1300_));
  NAND4_X1  g1108(.A1(new_n1257_), .A2(new_n1293_), .A3(new_n1294_), .A4(new_n1290_), .ZN(new_n1301_));
  NAND3_X1  g1109(.A1(new_n1299_), .A2(new_n1300_), .A3(new_n1301_), .ZN(new_n1302_));
  NAND3_X1  g1110(.A1(new_n1255_), .A2(new_n1296_), .A3(new_n1302_), .ZN(new_n1303_));
  NAND2_X1  g1111(.A1(new_n1117_), .A2(new_n1118_), .ZN(new_n1304_));
  INV_X1    g1112(.A(new_n1077_), .ZN(new_n1305_));
  OAI21_X1  g1113(.A(new_n1125_), .B1(new_n1304_), .B2(new_n1305_), .ZN(new_n1306_));
  INV_X1    g1114(.A(new_n1306_), .ZN(new_n1307_));
  NAND2_X1  g1115(.A1(new_n1303_), .A2(new_n1307_), .ZN(new_n1308_));
  NOR2_X1   g1116(.A1(new_n302_), .A2(new_n957_), .ZN(new_n1309_));
  INV_X1    g1117(.A(new_n1309_), .ZN(new_n1310_));
  NAND4_X1  g1118(.A1(new_n1306_), .A2(new_n1302_), .A3(new_n1255_), .A4(new_n1296_), .ZN(new_n1311_));
  AND3_X1   g1119(.A1(new_n1308_), .A2(new_n1310_), .A3(new_n1311_), .ZN(new_n1312_));
  AOI21_X1  g1120(.A(new_n1310_), .B1(new_n1308_), .B2(new_n1311_), .ZN(new_n1313_));
  NOR2_X1   g1121(.A1(new_n1312_), .A2(new_n1313_), .ZN(new_n1314_));
  AND3_X1   g1122(.A1(new_n1299_), .A2(new_n1300_), .A3(new_n1301_), .ZN(new_n1315_));
  AOI21_X1  g1123(.A(new_n1300_), .B1(new_n1299_), .B2(new_n1301_), .ZN(new_n1316_));
  NOR2_X1   g1124(.A1(new_n1315_), .A2(new_n1316_), .ZN(new_n1317_));
  AOI21_X1  g1125(.A(new_n1306_), .B1(new_n1317_), .B2(new_n1255_), .ZN(new_n1318_));
  AND4_X1   g1126(.A1(new_n1306_), .A2(new_n1302_), .A3(new_n1296_), .A4(new_n1255_), .ZN(new_n1319_));
  OAI21_X1  g1127(.A(new_n1310_), .B1(new_n1318_), .B2(new_n1319_), .ZN(new_n1320_));
  INV_X1    g1128(.A(KEYINPUT58), .ZN(new_n1321_));
  NAND2_X1  g1129(.A1(new_n1320_), .A2(new_n1321_), .ZN(new_n1322_));
  NAND2_X1  g1130(.A1(new_n1129_), .A2(new_n1128_), .ZN(new_n1323_));
  NAND3_X1  g1131(.A1(new_n1314_), .A2(new_n1322_), .A3(new_n1323_), .ZN(new_n1324_));
  NOR2_X1   g1132(.A1(new_n648_), .A2(new_n356_), .ZN(new_n1325_));
  INV_X1    g1133(.A(new_n1325_), .ZN(new_n1326_));
  AOI21_X1  g1134(.A(new_n1309_), .B1(new_n1308_), .B2(new_n1311_), .ZN(new_n1327_));
  OAI21_X1  g1135(.A(new_n1323_), .B1(new_n1327_), .B2(KEYINPUT58), .ZN(new_n1328_));
  OAI21_X1  g1136(.A(new_n1309_), .B1(new_n1318_), .B2(new_n1319_), .ZN(new_n1329_));
  NAND3_X1  g1137(.A1(new_n1308_), .A2(new_n1310_), .A3(new_n1311_), .ZN(new_n1330_));
  NAND2_X1  g1138(.A1(new_n1329_), .A2(new_n1330_), .ZN(new_n1331_));
  NAND2_X1  g1139(.A1(new_n1328_), .A2(new_n1331_), .ZN(new_n1332_));
  AND3_X1   g1140(.A1(new_n1324_), .A2(new_n1326_), .A3(new_n1332_), .ZN(new_n1333_));
  AOI21_X1  g1141(.A(new_n1326_), .B1(new_n1324_), .B2(new_n1332_), .ZN(new_n1334_));
  OAI21_X1  g1142(.A(new_n1253_), .B1(new_n1333_), .B2(new_n1334_), .ZN(new_n1335_));
  NOR2_X1   g1143(.A1(new_n539_), .A2(new_n867_), .ZN(new_n1336_));
  INV_X1    g1144(.A(new_n1336_), .ZN(new_n1337_));
  AND2_X1   g1145(.A1(new_n1328_), .A2(new_n1331_), .ZN(new_n1338_));
  NOR2_X1   g1146(.A1(new_n1328_), .A2(new_n1331_), .ZN(new_n1339_));
  OAI21_X1  g1147(.A(new_n1325_), .B1(new_n1338_), .B2(new_n1339_), .ZN(new_n1340_));
  NAND3_X1  g1148(.A1(new_n1324_), .A2(new_n1326_), .A3(new_n1332_), .ZN(new_n1341_));
  AND2_X1   g1149(.A1(new_n1245_), .A2(new_n1252_), .ZN(new_n1342_));
  NAND3_X1  g1150(.A1(new_n1340_), .A2(new_n1341_), .A3(new_n1342_), .ZN(new_n1343_));
  NAND3_X1  g1151(.A1(new_n1335_), .A2(new_n1337_), .A3(new_n1343_), .ZN(new_n1344_));
  AOI21_X1  g1152(.A(new_n1337_), .B1(new_n1335_), .B2(new_n1343_), .ZN(new_n1345_));
  INV_X1    g1153(.A(KEYINPUT59), .ZN(new_n1346_));
  OAI21_X1  g1154(.A(new_n1344_), .B1(new_n1345_), .B2(new_n1346_), .ZN(new_n1347_));
  AOI211_X1 g1155(.A(KEYINPUT59), .B(new_n1337_), .C1(new_n1335_), .C2(new_n1343_), .ZN(new_n1348_));
  OAI21_X1  g1156(.A(new_n1248_), .B1(new_n1347_), .B2(new_n1348_), .ZN(new_n1349_));
  NAND2_X1  g1157(.A1(new_n1335_), .A2(new_n1343_), .ZN(new_n1350_));
  NAND2_X1  g1158(.A1(new_n1350_), .A2(new_n1336_), .ZN(new_n1351_));
  NAND3_X1  g1159(.A1(new_n1351_), .A2(new_n1247_), .A3(new_n1344_), .ZN(new_n1352_));
  NAND2_X1  g1160(.A1(new_n1349_), .A2(new_n1352_), .ZN(new_n1353_));
  NOR2_X1   g1161(.A1(new_n455_), .A2(new_n616_), .ZN(new_n1354_));
  NAND2_X1  g1162(.A1(new_n1353_), .A2(new_n1354_), .ZN(new_n1355_));
  INV_X1    g1163(.A(KEYINPUT60), .ZN(new_n1356_));
  INV_X1    g1164(.A(new_n1354_), .ZN(new_n1357_));
  NAND3_X1  g1165(.A1(new_n1349_), .A2(new_n1357_), .A3(new_n1352_), .ZN(new_n1358_));
  NAND3_X1  g1166(.A1(new_n1355_), .A2(new_n1356_), .A3(new_n1358_), .ZN(new_n1359_));
  AOI21_X1  g1167(.A(new_n1161_), .B1(new_n1157_), .B2(new_n1156_), .ZN(new_n1360_));
  NAND3_X1  g1168(.A1(new_n1353_), .A2(KEYINPUT60), .A3(new_n1354_), .ZN(new_n1361_));
  NAND3_X1  g1169(.A1(new_n1359_), .A2(new_n1360_), .A3(new_n1361_), .ZN(new_n1362_));
  NOR2_X1   g1170(.A1(new_n312_), .A2(new_n774_), .ZN(new_n1363_));
  INV_X1    g1171(.A(new_n1360_), .ZN(new_n1364_));
  NAND3_X1  g1172(.A1(new_n1364_), .A2(new_n1355_), .A3(new_n1358_), .ZN(new_n1365_));
  AND3_X1   g1173(.A1(new_n1362_), .A2(new_n1363_), .A3(new_n1365_), .ZN(new_n1366_));
  AOI21_X1  g1174(.A(new_n1363_), .B1(new_n1362_), .B2(new_n1365_), .ZN(new_n1367_));
  NOR2_X1   g1175(.A1(new_n1366_), .A2(new_n1367_), .ZN(new_n1368_));
  NOR2_X1   g1176(.A1(new_n1024_), .A2(new_n1164_), .ZN(new_n1369_));
  NAND2_X1  g1177(.A1(new_n1163_), .A2(new_n1168_), .ZN(new_n1370_));
  NOR2_X1   g1178(.A1(new_n1369_), .A2(new_n1370_), .ZN(new_n1371_));
  INV_X1    g1179(.A(new_n1371_), .ZN(new_n1372_));
  NAND2_X1  g1180(.A1(new_n1187_), .A2(new_n1372_), .ZN(new_n1373_));
  NAND2_X1  g1181(.A1(new_n1368_), .A2(new_n1373_), .ZN(new_n1374_));
  NOR2_X1   g1182(.A1(new_n318_), .A2(new_n765_), .ZN(new_n1375_));
  INV_X1    g1183(.A(new_n1375_), .ZN(new_n1376_));
  OAI211_X1 g1184(.A(new_n1187_), .B(new_n1372_), .C1(new_n1366_), .C2(new_n1367_), .ZN(new_n1377_));
  AND3_X1   g1185(.A1(new_n1374_), .A2(new_n1376_), .A3(new_n1377_), .ZN(new_n1378_));
  AOI21_X1  g1186(.A(new_n1376_), .B1(new_n1374_), .B2(new_n1377_), .ZN(new_n1379_));
  OAI21_X1  g1187(.A(new_n1243_), .B1(new_n1378_), .B2(new_n1379_), .ZN(new_n1380_));
  INV_X1    g1188(.A(new_n1377_), .ZN(new_n1381_));
  AOI21_X1  g1189(.A(new_n1371_), .B1(new_n1184_), .B2(new_n1186_), .ZN(new_n1382_));
  NOR3_X1   g1190(.A1(new_n1382_), .A2(new_n1367_), .A3(new_n1366_), .ZN(new_n1383_));
  OAI21_X1  g1191(.A(new_n1375_), .B1(new_n1381_), .B2(new_n1383_), .ZN(new_n1384_));
  NAND3_X1  g1192(.A1(new_n1374_), .A2(new_n1376_), .A3(new_n1377_), .ZN(new_n1385_));
  NAND3_X1  g1193(.A1(new_n1384_), .A2(new_n1385_), .A3(new_n1242_), .ZN(new_n1386_));
  NOR2_X1   g1194(.A1(new_n214_), .A2(new_n1055_), .ZN(new_n1387_));
  AND3_X1   g1195(.A1(new_n1380_), .A2(new_n1386_), .A3(new_n1387_), .ZN(new_n1388_));
  XNOR2_X1  g1196(.A(new_n1387_), .B(KEYINPUT61), .ZN(new_n1389_));
  INV_X1    g1197(.A(new_n1389_), .ZN(new_n1390_));
  AOI21_X1  g1198(.A(new_n1390_), .B1(new_n1380_), .B2(new_n1386_), .ZN(new_n1391_));
  OAI21_X1  g1199(.A(new_n1241_), .B1(new_n1388_), .B2(new_n1391_), .ZN(new_n1392_));
  AND3_X1   g1200(.A1(new_n1384_), .A2(new_n1385_), .A3(new_n1242_), .ZN(new_n1393_));
  AOI21_X1  g1201(.A(new_n1242_), .B1(new_n1384_), .B2(new_n1385_), .ZN(new_n1394_));
  OAI21_X1  g1202(.A(new_n1389_), .B1(new_n1393_), .B2(new_n1394_), .ZN(new_n1395_));
  NAND3_X1  g1203(.A1(new_n1380_), .A2(new_n1386_), .A3(new_n1390_), .ZN(new_n1396_));
  NAND4_X1  g1204(.A1(new_n1395_), .A2(new_n1208_), .A3(new_n1240_), .A4(new_n1396_), .ZN(new_n1397_));
  NAND2_X1  g1205(.A1(new_n1392_), .A2(new_n1397_), .ZN(new_n1398_));
  NOR2_X1   g1206(.A1(new_n213_), .A2(new_n1215_), .ZN(new_n1399_));
  NAND2_X1  g1207(.A1(new_n1398_), .A2(new_n1399_), .ZN(new_n1400_));
  INV_X1    g1208(.A(new_n1399_), .ZN(new_n1401_));
  NAND3_X1  g1209(.A1(new_n1392_), .A2(new_n1401_), .A3(new_n1397_), .ZN(new_n1402_));
  AND2_X1   g1210(.A1(new_n1400_), .A2(new_n1402_), .ZN(new_n1403_));
  OR2_X1    g1211(.A1(new_n1236_), .A2(new_n1403_), .ZN(new_n1404_));
  INV_X1    g1212(.A(G494gat), .ZN(new_n1405_));
  NOR2_X1   g1213(.A1(new_n196_), .A2(new_n1405_), .ZN(new_n1406_));
  INV_X1    g1214(.A(new_n1406_), .ZN(new_n1407_));
  NAND3_X1  g1215(.A1(new_n1236_), .A2(new_n1400_), .A3(new_n1402_), .ZN(new_n1408_));
  NAND3_X1  g1216(.A1(new_n1404_), .A2(new_n1407_), .A3(new_n1408_), .ZN(new_n1409_));
  INV_X1    g1217(.A(new_n1409_), .ZN(new_n1410_));
  AOI21_X1  g1218(.A(new_n1407_), .B1(new_n1404_), .B2(new_n1408_), .ZN(new_n1411_));
  OAI211_X1 g1219(.A(new_n1232_), .B(new_n1227_), .C1(new_n1410_), .C2(new_n1411_), .ZN(new_n1412_));
  NAND3_X1  g1220(.A1(new_n1224_), .A2(new_n1227_), .A3(new_n1230_), .ZN(new_n1413_));
  INV_X1    g1221(.A(new_n1411_), .ZN(new_n1414_));
  NAND4_X1  g1222(.A1(new_n1413_), .A2(new_n1224_), .A3(new_n1414_), .A4(new_n1409_), .ZN(new_n1415_));
  NAND2_X1  g1223(.A1(new_n1412_), .A2(new_n1415_), .ZN(new_n1416_));
  INV_X1    g1224(.A(G511gat), .ZN(new_n1417_));
  NOR2_X1   g1225(.A1(new_n193_), .A2(new_n1417_), .ZN(new_n1418_));
  INV_X1    g1226(.A(new_n1418_), .ZN(new_n1419_));
  XNOR2_X1  g1227(.A(new_n1416_), .B(new_n1419_), .ZN(G5971gat));
  AND4_X1   g1228(.A1(new_n1227_), .A2(new_n1232_), .A3(new_n1409_), .A4(new_n1414_), .ZN(new_n1421_));
  AOI21_X1  g1229(.A(new_n1421_), .B1(new_n1416_), .B2(new_n1419_), .ZN(new_n1422_));
  NAND2_X1  g1230(.A1(G52gat), .A2(G477gat), .ZN(new_n1423_));
  NAND2_X1  g1231(.A1(new_n1362_), .A2(new_n1365_), .ZN(new_n1424_));
  INV_X1    g1232(.A(new_n1363_), .ZN(new_n1425_));
  NAND2_X1  g1233(.A1(new_n1424_), .A2(new_n1425_), .ZN(new_n1426_));
  NAND3_X1  g1234(.A1(new_n1359_), .A2(new_n1364_), .A3(new_n1361_), .ZN(new_n1427_));
  NAND2_X1  g1235(.A1(new_n1317_), .A2(new_n1306_), .ZN(new_n1428_));
  NAND2_X1  g1236(.A1(new_n1289_), .A2(new_n1257_), .ZN(new_n1429_));
  INV_X1    g1237(.A(KEYINPUT66), .ZN(new_n1430_));
  NAND2_X1  g1238(.A1(G239gat), .A2(G290gat), .ZN(new_n1431_));
  AOI21_X1  g1239(.A(new_n1431_), .B1(G256gat), .B2(G273gat), .ZN(new_n1432_));
  NAND2_X1  g1240(.A1(new_n1432_), .A2(new_n1261_), .ZN(new_n1433_));
  NAND2_X1  g1241(.A1(G256gat), .A2(G273gat), .ZN(new_n1434_));
  OAI21_X1  g1242(.A(new_n1259_), .B1(new_n1262_), .B2(new_n1434_), .ZN(new_n1435_));
  OAI21_X1  g1243(.A(new_n1433_), .B1(new_n1432_), .B2(new_n1435_), .ZN(new_n1436_));
  INV_X1    g1244(.A(G222gat), .ZN(new_n1437_));
  NOR2_X1   g1245(.A1(new_n1437_), .A2(new_n245_), .ZN(new_n1438_));
  NAND2_X1  g1246(.A1(new_n1436_), .A2(new_n1438_), .ZN(new_n1439_));
  INV_X1    g1247(.A(new_n1438_), .ZN(new_n1440_));
  OAI211_X1 g1248(.A(new_n1433_), .B(new_n1440_), .C1(new_n1432_), .C2(new_n1435_), .ZN(new_n1441_));
  NAND2_X1  g1249(.A1(new_n1439_), .A2(new_n1441_), .ZN(new_n1442_));
  INV_X1    g1250(.A(new_n1442_), .ZN(new_n1443_));
  NAND2_X1  g1251(.A1(new_n1283_), .A2(new_n1268_), .ZN(new_n1444_));
  NAND2_X1  g1252(.A1(new_n1444_), .A2(KEYINPUT65), .ZN(new_n1445_));
  INV_X1    g1253(.A(new_n1276_), .ZN(new_n1446_));
  AOI21_X1  g1254(.A(new_n1267_), .B1(new_n1266_), .B2(new_n1271_), .ZN(new_n1447_));
  INV_X1    g1255(.A(KEYINPUT65), .ZN(new_n1448_));
  AOI21_X1  g1256(.A(new_n1446_), .B1(new_n1447_), .B2(new_n1448_), .ZN(new_n1449_));
  AOI21_X1  g1257(.A(new_n1443_), .B1(new_n1445_), .B2(new_n1449_), .ZN(new_n1450_));
  NOR2_X1   g1258(.A1(new_n1438_), .A2(KEYINPUT64), .ZN(new_n1451_));
  NAND2_X1  g1259(.A1(new_n1436_), .A2(new_n1451_), .ZN(new_n1452_));
  INV_X1    g1260(.A(new_n1260_), .ZN(new_n1453_));
  OAI211_X1 g1261(.A(new_n1452_), .B(new_n1276_), .C1(new_n1267_), .C2(new_n1453_), .ZN(new_n1454_));
  INV_X1    g1262(.A(KEYINPUT64), .ZN(new_n1455_));
  AOI21_X1  g1263(.A(new_n1455_), .B1(new_n1439_), .B2(new_n1441_), .ZN(new_n1456_));
  NOR2_X1   g1264(.A1(new_n1454_), .A2(new_n1456_), .ZN(new_n1457_));
  OAI21_X1  g1265(.A(new_n1430_), .B1(new_n1450_), .B2(new_n1457_), .ZN(new_n1458_));
  NAND3_X1  g1266(.A1(new_n1283_), .A2(new_n1448_), .A3(new_n1268_), .ZN(new_n1459_));
  NAND2_X1  g1267(.A1(new_n1459_), .A2(new_n1276_), .ZN(new_n1460_));
  NOR2_X1   g1268(.A1(new_n1447_), .A2(new_n1448_), .ZN(new_n1461_));
  OAI21_X1  g1269(.A(new_n1442_), .B1(new_n1460_), .B2(new_n1461_), .ZN(new_n1462_));
  OR2_X1    g1270(.A1(new_n1454_), .A2(new_n1456_), .ZN(new_n1463_));
  NAND3_X1  g1271(.A1(new_n1462_), .A2(KEYINPUT66), .A3(new_n1463_), .ZN(new_n1464_));
  NOR2_X1   g1272(.A1(new_n942_), .A2(new_n232_), .ZN(new_n1465_));
  NAND3_X1  g1273(.A1(new_n1458_), .A2(new_n1464_), .A3(new_n1465_), .ZN(new_n1466_));
  AOI22_X1  g1274(.A1(new_n1286_), .A2(new_n1282_), .B1(new_n1279_), .B2(new_n1278_), .ZN(new_n1467_));
  NOR2_X1   g1275(.A1(new_n1450_), .A2(new_n1457_), .ZN(new_n1468_));
  INV_X1    g1276(.A(new_n1465_), .ZN(new_n1469_));
  AOI21_X1  g1277(.A(new_n1467_), .B1(new_n1468_), .B2(new_n1469_), .ZN(new_n1470_));
  NAND2_X1  g1278(.A1(new_n1466_), .A2(new_n1470_), .ZN(new_n1471_));
  NOR2_X1   g1279(.A1(new_n1092_), .A2(new_n261_), .ZN(new_n1472_));
  OAI21_X1  g1280(.A(new_n1465_), .B1(new_n1450_), .B2(new_n1457_), .ZN(new_n1473_));
  NAND3_X1  g1281(.A1(new_n1462_), .A2(new_n1469_), .A3(new_n1463_), .ZN(new_n1474_));
  NAND2_X1  g1282(.A1(new_n1473_), .A2(new_n1474_), .ZN(new_n1475_));
  NAND2_X1  g1283(.A1(new_n1475_), .A2(new_n1467_), .ZN(new_n1476_));
  AND3_X1   g1284(.A1(new_n1471_), .A2(new_n1472_), .A3(new_n1476_), .ZN(new_n1477_));
  AOI21_X1  g1285(.A(new_n1472_), .B1(new_n1471_), .B2(new_n1476_), .ZN(new_n1478_));
  OAI211_X1 g1286(.A(new_n1302_), .B(new_n1429_), .C1(new_n1477_), .C2(new_n1478_), .ZN(new_n1479_));
  NOR2_X1   g1287(.A1(new_n302_), .A2(new_n946_), .ZN(new_n1480_));
  INV_X1    g1288(.A(new_n1480_), .ZN(new_n1481_));
  NAND2_X1  g1289(.A1(new_n1471_), .A2(new_n1476_), .ZN(new_n1482_));
  INV_X1    g1290(.A(new_n1472_), .ZN(new_n1483_));
  NAND2_X1  g1291(.A1(new_n1482_), .A2(new_n1483_), .ZN(new_n1484_));
  NAND2_X1  g1292(.A1(new_n1302_), .A2(new_n1429_), .ZN(new_n1485_));
  AOI22_X1  g1293(.A1(new_n1466_), .A2(new_n1470_), .B1(new_n1475_), .B2(new_n1467_), .ZN(new_n1486_));
  NAND2_X1  g1294(.A1(new_n1486_), .A2(new_n1472_), .ZN(new_n1487_));
  NAND3_X1  g1295(.A1(new_n1484_), .A2(new_n1485_), .A3(new_n1487_), .ZN(new_n1488_));
  AND3_X1   g1296(.A1(new_n1479_), .A2(new_n1481_), .A3(new_n1488_), .ZN(new_n1489_));
  AOI21_X1  g1297(.A(new_n1481_), .B1(new_n1479_), .B2(new_n1488_), .ZN(new_n1490_));
  OAI211_X1 g1298(.A(new_n1330_), .B(new_n1428_), .C1(new_n1489_), .C2(new_n1490_), .ZN(new_n1491_));
  NAND2_X1  g1299(.A1(new_n1330_), .A2(new_n1428_), .ZN(new_n1492_));
  NAND3_X1  g1300(.A1(new_n1479_), .A2(new_n1488_), .A3(new_n1481_), .ZN(new_n1493_));
  INV_X1    g1301(.A(new_n1488_), .ZN(new_n1494_));
  AOI21_X1  g1302(.A(new_n1485_), .B1(new_n1484_), .B2(new_n1487_), .ZN(new_n1495_));
  OAI21_X1  g1303(.A(new_n1480_), .B1(new_n1494_), .B2(new_n1495_), .ZN(new_n1496_));
  NAND3_X1  g1304(.A1(new_n1492_), .A2(new_n1493_), .A3(new_n1496_), .ZN(new_n1497_));
  NOR2_X1   g1305(.A1(new_n957_), .A2(new_n356_), .ZN(new_n1498_));
  INV_X1    g1306(.A(new_n1498_), .ZN(new_n1499_));
  AND3_X1   g1307(.A1(new_n1491_), .A2(new_n1497_), .A3(new_n1499_), .ZN(new_n1500_));
  AOI21_X1  g1308(.A(new_n1499_), .B1(new_n1491_), .B2(new_n1497_), .ZN(new_n1501_));
  NOR2_X1   g1309(.A1(new_n1500_), .A2(new_n1501_), .ZN(new_n1502_));
  NAND2_X1  g1310(.A1(new_n1314_), .A2(new_n1323_), .ZN(new_n1503_));
  NAND2_X1  g1311(.A1(new_n1341_), .A2(new_n1503_), .ZN(new_n1504_));
  NAND2_X1  g1312(.A1(new_n1502_), .A2(new_n1504_), .ZN(new_n1505_));
  OAI211_X1 g1313(.A(new_n1341_), .B(new_n1503_), .C1(new_n1500_), .C2(new_n1501_), .ZN(new_n1506_));
  NAND2_X1  g1314(.A1(new_n1505_), .A2(new_n1506_), .ZN(new_n1507_));
  NOR2_X1   g1315(.A1(new_n648_), .A2(new_n867_), .ZN(new_n1508_));
  NAND2_X1  g1316(.A1(new_n1507_), .A2(new_n1508_), .ZN(new_n1509_));
  INV_X1    g1317(.A(new_n1508_), .ZN(new_n1510_));
  NAND3_X1  g1318(.A1(new_n1505_), .A2(new_n1510_), .A3(new_n1506_), .ZN(new_n1511_));
  AOI21_X1  g1319(.A(new_n1336_), .B1(new_n1335_), .B2(new_n1343_), .ZN(new_n1512_));
  NAND3_X1  g1320(.A1(new_n1340_), .A2(new_n1341_), .A3(new_n1253_), .ZN(new_n1513_));
  INV_X1    g1321(.A(new_n1513_), .ZN(new_n1514_));
  OAI211_X1 g1322(.A(new_n1509_), .B(new_n1511_), .C1(new_n1512_), .C2(new_n1514_), .ZN(new_n1515_));
  AND3_X1   g1323(.A1(new_n1340_), .A2(new_n1341_), .A3(new_n1342_), .ZN(new_n1516_));
  AOI22_X1  g1324(.A1(new_n1340_), .A2(new_n1341_), .B1(new_n1149_), .B2(new_n1252_), .ZN(new_n1517_));
  OAI21_X1  g1325(.A(new_n1337_), .B1(new_n1516_), .B2(new_n1517_), .ZN(new_n1518_));
  AND3_X1   g1326(.A1(new_n1505_), .A2(new_n1510_), .A3(new_n1506_), .ZN(new_n1519_));
  AOI21_X1  g1327(.A(new_n1510_), .B1(new_n1505_), .B2(new_n1506_), .ZN(new_n1520_));
  OAI211_X1 g1328(.A(new_n1518_), .B(new_n1513_), .C1(new_n1519_), .C2(new_n1520_), .ZN(new_n1521_));
  NOR2_X1   g1329(.A1(new_n539_), .A2(new_n616_), .ZN(new_n1522_));
  INV_X1    g1330(.A(new_n1522_), .ZN(new_n1523_));
  NAND3_X1  g1331(.A1(new_n1515_), .A2(new_n1521_), .A3(new_n1523_), .ZN(new_n1524_));
  INV_X1    g1332(.A(new_n1524_), .ZN(new_n1525_));
  AOI21_X1  g1333(.A(new_n1523_), .B1(new_n1515_), .B2(new_n1521_), .ZN(new_n1526_));
  OR2_X1    g1334(.A1(new_n1525_), .A2(new_n1526_), .ZN(new_n1527_));
  NAND2_X1  g1335(.A1(new_n1351_), .A2(KEYINPUT59), .ZN(new_n1528_));
  NAND2_X1  g1336(.A1(new_n1345_), .A2(new_n1346_), .ZN(new_n1529_));
  NAND3_X1  g1337(.A1(new_n1528_), .A2(new_n1529_), .A3(new_n1344_), .ZN(new_n1530_));
  NAND2_X1  g1338(.A1(new_n1530_), .A2(new_n1247_), .ZN(new_n1531_));
  AOI21_X1  g1339(.A(new_n1354_), .B1(new_n1349_), .B2(new_n1352_), .ZN(new_n1532_));
  INV_X1    g1340(.A(KEYINPUT67), .ZN(new_n1533_));
  OAI21_X1  g1341(.A(new_n1531_), .B1(new_n1532_), .B2(new_n1533_), .ZN(new_n1534_));
  AOI211_X1 g1342(.A(KEYINPUT67), .B(new_n1354_), .C1(new_n1349_), .C2(new_n1352_), .ZN(new_n1535_));
  OAI21_X1  g1343(.A(new_n1527_), .B1(new_n1534_), .B2(new_n1535_), .ZN(new_n1536_));
  NOR2_X1   g1344(.A1(new_n455_), .A2(new_n774_), .ZN(new_n1537_));
  NOR2_X1   g1345(.A1(new_n1525_), .A2(new_n1526_), .ZN(new_n1538_));
  NAND2_X1  g1346(.A1(new_n1353_), .A2(new_n1357_), .ZN(new_n1539_));
  NAND3_X1  g1347(.A1(new_n1538_), .A2(new_n1539_), .A3(new_n1531_), .ZN(new_n1540_));
  NAND3_X1  g1348(.A1(new_n1536_), .A2(new_n1537_), .A3(new_n1540_), .ZN(new_n1541_));
  INV_X1    g1349(.A(new_n1541_), .ZN(new_n1542_));
  AOI21_X1  g1350(.A(new_n1537_), .B1(new_n1536_), .B2(new_n1540_), .ZN(new_n1543_));
  OAI211_X1 g1351(.A(new_n1426_), .B(new_n1427_), .C1(new_n1542_), .C2(new_n1543_), .ZN(new_n1544_));
  INV_X1    g1352(.A(new_n1537_), .ZN(new_n1545_));
  AND2_X1   g1353(.A1(new_n1530_), .A2(new_n1247_), .ZN(new_n1546_));
  AOI21_X1  g1354(.A(new_n1546_), .B1(new_n1539_), .B2(KEYINPUT67), .ZN(new_n1547_));
  INV_X1    g1355(.A(new_n1535_), .ZN(new_n1548_));
  AOI21_X1  g1356(.A(new_n1538_), .B1(new_n1547_), .B2(new_n1548_), .ZN(new_n1549_));
  INV_X1    g1357(.A(new_n1540_), .ZN(new_n1550_));
  OAI21_X1  g1358(.A(new_n1545_), .B1(new_n1549_), .B2(new_n1550_), .ZN(new_n1551_));
  INV_X1    g1359(.A(new_n1427_), .ZN(new_n1552_));
  OAI211_X1 g1360(.A(new_n1551_), .B(new_n1541_), .C1(new_n1367_), .C2(new_n1552_), .ZN(new_n1553_));
  NOR2_X1   g1361(.A1(new_n312_), .A2(new_n765_), .ZN(new_n1554_));
  NAND3_X1  g1362(.A1(new_n1544_), .A2(new_n1553_), .A3(new_n1554_), .ZN(new_n1555_));
  NAND2_X1  g1363(.A1(new_n1555_), .A2(KEYINPUT68), .ZN(new_n1556_));
  OAI21_X1  g1364(.A(new_n1374_), .B1(new_n1381_), .B2(new_n1375_), .ZN(new_n1557_));
  NAND2_X1  g1365(.A1(new_n1556_), .A2(new_n1557_), .ZN(new_n1558_));
  NAND2_X1  g1366(.A1(new_n1544_), .A2(new_n1553_), .ZN(new_n1559_));
  NAND2_X1  g1367(.A1(new_n1559_), .A2(new_n1554_), .ZN(new_n1560_));
  INV_X1    g1368(.A(new_n1554_), .ZN(new_n1561_));
  NAND3_X1  g1369(.A1(new_n1544_), .A2(new_n1553_), .A3(new_n1561_), .ZN(new_n1562_));
  NAND2_X1  g1370(.A1(new_n1560_), .A2(new_n1562_), .ZN(new_n1563_));
  NAND2_X1  g1371(.A1(new_n1558_), .A2(new_n1563_), .ZN(new_n1564_));
  NOR2_X1   g1372(.A1(new_n318_), .A2(new_n1055_), .ZN(new_n1565_));
  INV_X1    g1373(.A(new_n1565_), .ZN(new_n1566_));
  NAND4_X1  g1374(.A1(new_n1556_), .A2(new_n1557_), .A3(new_n1560_), .A4(new_n1562_), .ZN(new_n1567_));
  AND3_X1   g1375(.A1(new_n1564_), .A2(new_n1566_), .A3(new_n1567_), .ZN(new_n1568_));
  AOI21_X1  g1376(.A(new_n1566_), .B1(new_n1564_), .B2(new_n1567_), .ZN(new_n1569_));
  NAND2_X1  g1377(.A1(new_n1380_), .A2(new_n1389_), .ZN(new_n1570_));
  NAND2_X1  g1378(.A1(new_n1570_), .A2(new_n1386_), .ZN(new_n1571_));
  NOR3_X1   g1379(.A1(new_n1568_), .A2(new_n1569_), .A3(new_n1571_), .ZN(new_n1572_));
  INV_X1    g1380(.A(new_n1387_), .ZN(new_n1573_));
  OAI21_X1  g1381(.A(new_n1380_), .B1(new_n1393_), .B2(new_n1573_), .ZN(new_n1574_));
  NOR2_X1   g1382(.A1(new_n1558_), .A2(new_n1563_), .ZN(new_n1575_));
  AOI22_X1  g1383(.A1(new_n1556_), .A2(new_n1557_), .B1(new_n1560_), .B2(new_n1562_), .ZN(new_n1576_));
  OAI21_X1  g1384(.A(new_n1565_), .B1(new_n1575_), .B2(new_n1576_), .ZN(new_n1577_));
  NAND3_X1  g1385(.A1(new_n1564_), .A2(new_n1566_), .A3(new_n1567_), .ZN(new_n1578_));
  AOI21_X1  g1386(.A(new_n1574_), .B1(new_n1577_), .B2(new_n1578_), .ZN(new_n1579_));
  OAI21_X1  g1387(.A(new_n1423_), .B1(new_n1572_), .B2(new_n1579_), .ZN(new_n1580_));
  INV_X1    g1388(.A(new_n1574_), .ZN(new_n1581_));
  OAI21_X1  g1389(.A(new_n1581_), .B1(new_n1568_), .B2(new_n1569_), .ZN(new_n1582_));
  NAND4_X1  g1390(.A1(new_n1577_), .A2(new_n1386_), .A3(new_n1578_), .A4(new_n1570_), .ZN(new_n1583_));
  NAND4_X1  g1391(.A1(new_n1582_), .A2(new_n1583_), .A3(G52gat), .A4(G477gat), .ZN(new_n1584_));
  INV_X1    g1392(.A(new_n1396_), .ZN(new_n1585_));
  OAI21_X1  g1393(.A(new_n1241_), .B1(new_n1585_), .B2(new_n1391_), .ZN(new_n1586_));
  AOI22_X1  g1394(.A1(new_n1580_), .A2(new_n1584_), .B1(new_n1402_), .B2(new_n1586_), .ZN(new_n1587_));
  NAND2_X1  g1395(.A1(new_n1402_), .A2(KEYINPUT62), .ZN(new_n1588_));
  INV_X1    g1396(.A(KEYINPUT62), .ZN(new_n1589_));
  NAND4_X1  g1397(.A1(new_n1392_), .A2(new_n1397_), .A3(new_n1589_), .A4(new_n1401_), .ZN(new_n1590_));
  INV_X1    g1398(.A(KEYINPUT63), .ZN(new_n1591_));
  NAND2_X1  g1399(.A1(new_n1586_), .A2(new_n1591_), .ZN(new_n1592_));
  OAI211_X1 g1400(.A(new_n1241_), .B(KEYINPUT63), .C1(new_n1585_), .C2(new_n1391_), .ZN(new_n1593_));
  NAND2_X1  g1401(.A1(new_n1592_), .A2(new_n1593_), .ZN(new_n1594_));
  AND3_X1   g1402(.A1(new_n1588_), .A2(new_n1590_), .A3(new_n1594_), .ZN(new_n1595_));
  NAND2_X1  g1403(.A1(new_n1580_), .A2(new_n1584_), .ZN(new_n1596_));
  INV_X1    g1404(.A(new_n1596_), .ZN(new_n1597_));
  AOI21_X1  g1405(.A(new_n1587_), .B1(new_n1595_), .B2(new_n1597_), .ZN(new_n1598_));
  NOR2_X1   g1406(.A1(new_n213_), .A2(new_n1405_), .ZN(new_n1599_));
  NOR2_X1   g1407(.A1(new_n1598_), .A2(new_n1599_), .ZN(new_n1600_));
  NAND2_X1  g1408(.A1(new_n1402_), .A2(new_n1586_), .ZN(new_n1601_));
  NAND2_X1  g1409(.A1(new_n1596_), .A2(new_n1601_), .ZN(new_n1602_));
  NAND3_X1  g1410(.A1(new_n1588_), .A2(new_n1590_), .A3(new_n1594_), .ZN(new_n1603_));
  OAI211_X1 g1411(.A(new_n1602_), .B(new_n1599_), .C1(new_n1596_), .C2(new_n1603_), .ZN(new_n1604_));
  INV_X1    g1412(.A(new_n1604_), .ZN(new_n1605_));
  OAI211_X1 g1413(.A(new_n1408_), .B(new_n1409_), .C1(new_n1600_), .C2(new_n1605_), .ZN(new_n1606_));
  NOR2_X1   g1414(.A1(new_n1236_), .A2(new_n1403_), .ZN(new_n1607_));
  OAI21_X1  g1415(.A(new_n1408_), .B1(new_n1607_), .B2(new_n1406_), .ZN(new_n1608_));
  OAI21_X1  g1416(.A(new_n1602_), .B1(new_n1596_), .B2(new_n1603_), .ZN(new_n1609_));
  INV_X1    g1417(.A(new_n1599_), .ZN(new_n1610_));
  NAND2_X1  g1418(.A1(new_n1609_), .A2(new_n1610_), .ZN(new_n1611_));
  NAND3_X1  g1419(.A1(new_n1608_), .A2(new_n1611_), .A3(new_n1604_), .ZN(new_n1612_));
  NAND2_X1  g1420(.A1(new_n1606_), .A2(new_n1612_), .ZN(new_n1613_));
  NAND3_X1  g1421(.A1(new_n1613_), .A2(G18gat), .A3(G511gat), .ZN(new_n1614_));
  NAND2_X1  g1422(.A1(G18gat), .A2(G511gat), .ZN(new_n1615_));
  NAND3_X1  g1423(.A1(new_n1606_), .A2(new_n1615_), .A3(new_n1612_), .ZN(new_n1616_));
  NAND2_X1  g1424(.A1(new_n1614_), .A2(new_n1616_), .ZN(new_n1617_));
  NOR2_X1   g1425(.A1(new_n1422_), .A2(new_n1617_), .ZN(new_n1618_));
  INV_X1    g1426(.A(new_n1618_), .ZN(new_n1619_));
  NAND2_X1  g1427(.A1(new_n1422_), .A2(new_n1617_), .ZN(new_n1620_));
  NAND2_X1  g1428(.A1(new_n1619_), .A2(new_n1620_), .ZN(new_n1621_));
  INV_X1    g1429(.A(G528gat), .ZN(new_n1622_));
  NOR2_X1   g1430(.A1(new_n193_), .A2(new_n1622_), .ZN(new_n1623_));
  XNOR2_X1  g1431(.A(new_n1621_), .B(new_n1623_), .ZN(G6123gat));
  OAI21_X1  g1432(.A(KEYINPUT69), .B1(new_n1600_), .B2(new_n1605_), .ZN(new_n1625_));
  INV_X1    g1433(.A(KEYINPUT69), .ZN(new_n1626_));
  NAND3_X1  g1434(.A1(new_n1611_), .A2(new_n1626_), .A3(new_n1604_), .ZN(new_n1627_));
  NAND3_X1  g1435(.A1(new_n1625_), .A2(new_n1627_), .A3(new_n1608_), .ZN(new_n1628_));
  NAND2_X1  g1436(.A1(new_n1616_), .A2(new_n1628_), .ZN(new_n1629_));
  NAND3_X1  g1437(.A1(new_n1557_), .A2(new_n1560_), .A3(new_n1562_), .ZN(new_n1630_));
  NAND2_X1  g1438(.A1(new_n1578_), .A2(new_n1630_), .ZN(new_n1631_));
  INV_X1    g1439(.A(new_n1553_), .ZN(new_n1632_));
  AOI21_X1  g1440(.A(new_n1632_), .B1(new_n1561_), .B2(new_n1544_), .ZN(new_n1633_));
  AOI21_X1  g1441(.A(new_n1527_), .B1(new_n1547_), .B2(new_n1548_), .ZN(new_n1634_));
  INV_X1    g1442(.A(new_n1634_), .ZN(new_n1635_));
  NAND2_X1  g1443(.A1(new_n1551_), .A2(new_n1635_), .ZN(new_n1636_));
  INV_X1    g1444(.A(KEYINPUT72), .ZN(new_n1637_));
  NOR2_X1   g1445(.A1(new_n1519_), .A2(new_n1520_), .ZN(new_n1638_));
  NAND2_X1  g1446(.A1(new_n1518_), .A2(new_n1513_), .ZN(new_n1639_));
  NOR2_X1   g1447(.A1(new_n1638_), .A2(new_n1639_), .ZN(new_n1640_));
  OAI21_X1  g1448(.A(new_n1515_), .B1(new_n1640_), .B2(new_n1522_), .ZN(new_n1641_));
  NAND2_X1  g1449(.A1(G154gat), .A2(G392gat), .ZN(new_n1642_));
  AND3_X1   g1450(.A1(new_n1492_), .A2(new_n1493_), .A3(new_n1496_), .ZN(new_n1643_));
  AOI21_X1  g1451(.A(new_n1643_), .B1(new_n1499_), .B2(new_n1491_), .ZN(new_n1644_));
  AOI21_X1  g1452(.A(new_n1494_), .B1(new_n1481_), .B2(new_n1479_), .ZN(new_n1645_));
  INV_X1    g1453(.A(new_n1467_), .ZN(new_n1646_));
  AOI22_X1  g1454(.A1(new_n1482_), .A2(new_n1483_), .B1(new_n1646_), .B2(new_n1475_), .ZN(new_n1647_));
  NOR2_X1   g1455(.A1(new_n942_), .A2(new_n261_), .ZN(new_n1648_));
  INV_X1    g1456(.A(new_n1648_), .ZN(new_n1649_));
  NAND3_X1  g1457(.A1(new_n1458_), .A2(new_n1464_), .A3(new_n1469_), .ZN(new_n1650_));
  OAI21_X1  g1458(.A(new_n1276_), .B1(new_n1453_), .B2(new_n1267_), .ZN(new_n1651_));
  NAND2_X1  g1459(.A1(new_n1443_), .A2(new_n1651_), .ZN(new_n1652_));
  NAND2_X1  g1460(.A1(new_n1650_), .A2(new_n1652_), .ZN(new_n1653_));
  AND3_X1   g1461(.A1(new_n1261_), .A2(new_n1262_), .A3(new_n1434_), .ZN(new_n1654_));
  OAI22_X1  g1462(.A1(new_n1654_), .A2(new_n1438_), .B1(new_n1435_), .B2(new_n1432_), .ZN(new_n1655_));
  NAND3_X1  g1463(.A1(new_n1264_), .A2(G256gat), .A3(G290gat), .ZN(new_n1656_));
  INV_X1    g1464(.A(G239gat), .ZN(new_n1657_));
  NOR2_X1   g1465(.A1(new_n1657_), .A2(new_n245_), .ZN(new_n1658_));
  XNOR2_X1  g1466(.A(new_n1656_), .B(new_n1658_), .ZN(new_n1659_));
  NOR2_X1   g1467(.A1(new_n1655_), .A2(new_n1659_), .ZN(new_n1660_));
  INV_X1    g1468(.A(KEYINPUT70), .ZN(new_n1661_));
  OR3_X1    g1469(.A1(new_n1435_), .A2(new_n1432_), .A3(new_n1661_), .ZN(new_n1662_));
  OAI21_X1  g1470(.A(new_n1661_), .B1(new_n1435_), .B2(new_n1432_), .ZN(new_n1663_));
  NAND3_X1  g1471(.A1(new_n1441_), .A2(new_n1662_), .A3(new_n1663_), .ZN(new_n1664_));
  AOI21_X1  g1472(.A(new_n1660_), .B1(new_n1664_), .B2(new_n1659_), .ZN(new_n1665_));
  NOR2_X1   g1473(.A1(new_n1437_), .A2(new_n232_), .ZN(new_n1666_));
  INV_X1    g1474(.A(new_n1666_), .ZN(new_n1667_));
  INV_X1    g1475(.A(new_n1659_), .ZN(new_n1668_));
  OAI21_X1  g1476(.A(new_n1667_), .B1(new_n1668_), .B2(new_n1655_), .ZN(new_n1669_));
  INV_X1    g1477(.A(new_n1669_), .ZN(new_n1670_));
  NAND2_X1  g1478(.A1(new_n1664_), .A2(new_n1668_), .ZN(new_n1671_));
  AOI22_X1  g1479(.A1(new_n1665_), .A2(new_n1666_), .B1(new_n1670_), .B2(new_n1671_), .ZN(new_n1672_));
  NAND2_X1  g1480(.A1(new_n1653_), .A2(new_n1672_), .ZN(new_n1673_));
  INV_X1    g1481(.A(new_n1672_), .ZN(new_n1674_));
  OAI211_X1 g1482(.A(new_n1652_), .B(new_n1674_), .C1(new_n1468_), .C2(new_n1465_), .ZN(new_n1675_));
  AOI21_X1  g1483(.A(new_n1649_), .B1(new_n1673_), .B2(new_n1675_), .ZN(new_n1676_));
  AOI21_X1  g1484(.A(new_n1674_), .B1(new_n1650_), .B2(new_n1652_), .ZN(new_n1677_));
  INV_X1    g1485(.A(new_n1675_), .ZN(new_n1678_));
  NOR3_X1   g1486(.A1(new_n1677_), .A2(new_n1648_), .A3(new_n1678_), .ZN(new_n1679_));
  OAI21_X1  g1487(.A(new_n1647_), .B1(new_n1676_), .B2(new_n1679_), .ZN(new_n1680_));
  NOR2_X1   g1488(.A1(new_n302_), .A2(new_n1092_), .ZN(new_n1681_));
  INV_X1    g1489(.A(new_n1681_), .ZN(new_n1682_));
  NAND3_X1  g1490(.A1(new_n1673_), .A2(new_n1649_), .A3(new_n1675_), .ZN(new_n1683_));
  NAND2_X1  g1491(.A1(new_n1475_), .A2(new_n1646_), .ZN(new_n1684_));
  OAI21_X1  g1492(.A(new_n1684_), .B1(new_n1486_), .B2(new_n1472_), .ZN(new_n1685_));
  OAI21_X1  g1493(.A(new_n1648_), .B1(new_n1677_), .B2(new_n1678_), .ZN(new_n1686_));
  NAND3_X1  g1494(.A1(new_n1683_), .A2(new_n1685_), .A3(new_n1686_), .ZN(new_n1687_));
  AND3_X1   g1495(.A1(new_n1680_), .A2(new_n1682_), .A3(new_n1687_), .ZN(new_n1688_));
  AOI21_X1  g1496(.A(new_n1682_), .B1(new_n1680_), .B2(new_n1687_), .ZN(new_n1689_));
  OAI21_X1  g1497(.A(new_n1645_), .B1(new_n1688_), .B2(new_n1689_), .ZN(new_n1690_));
  NAND2_X1  g1498(.A1(new_n1680_), .A2(new_n1687_), .ZN(new_n1691_));
  NAND2_X1  g1499(.A1(new_n1691_), .A2(new_n1681_), .ZN(new_n1692_));
  NAND2_X1  g1500(.A1(new_n1493_), .A2(new_n1488_), .ZN(new_n1693_));
  NAND3_X1  g1501(.A1(new_n1680_), .A2(new_n1682_), .A3(new_n1687_), .ZN(new_n1694_));
  NAND3_X1  g1502(.A1(new_n1692_), .A2(new_n1693_), .A3(new_n1694_), .ZN(new_n1695_));
  NOR2_X1   g1503(.A1(new_n946_), .A2(new_n356_), .ZN(new_n1696_));
  INV_X1    g1504(.A(new_n1696_), .ZN(new_n1697_));
  AND3_X1   g1505(.A1(new_n1690_), .A2(new_n1695_), .A3(new_n1697_), .ZN(new_n1698_));
  AOI21_X1  g1506(.A(new_n1697_), .B1(new_n1690_), .B2(new_n1695_), .ZN(new_n1699_));
  OAI21_X1  g1507(.A(new_n1644_), .B1(new_n1698_), .B2(new_n1699_), .ZN(new_n1700_));
  NOR3_X1   g1508(.A1(new_n1688_), .A2(new_n1645_), .A3(new_n1689_), .ZN(new_n1701_));
  AOI21_X1  g1509(.A(new_n1693_), .B1(new_n1692_), .B2(new_n1694_), .ZN(new_n1702_));
  OAI21_X1  g1510(.A(new_n1696_), .B1(new_n1701_), .B2(new_n1702_), .ZN(new_n1703_));
  AOI21_X1  g1511(.A(new_n1492_), .B1(new_n1493_), .B2(new_n1496_), .ZN(new_n1704_));
  OAI21_X1  g1512(.A(new_n1497_), .B1(new_n1704_), .B2(new_n1498_), .ZN(new_n1705_));
  NAND3_X1  g1513(.A1(new_n1690_), .A2(new_n1695_), .A3(new_n1697_), .ZN(new_n1706_));
  NAND3_X1  g1514(.A1(new_n1703_), .A2(new_n1705_), .A3(new_n1706_), .ZN(new_n1707_));
  AOI21_X1  g1515(.A(new_n1642_), .B1(new_n1700_), .B2(new_n1707_), .ZN(new_n1708_));
  INV_X1    g1516(.A(new_n1708_), .ZN(new_n1709_));
  INV_X1    g1517(.A(new_n1506_), .ZN(new_n1710_));
  OAI21_X1  g1518(.A(new_n1505_), .B1(new_n1710_), .B2(new_n1508_), .ZN(new_n1711_));
  NAND3_X1  g1519(.A1(new_n1700_), .A2(new_n1707_), .A3(new_n1642_), .ZN(new_n1712_));
  NAND3_X1  g1520(.A1(new_n1709_), .A2(new_n1711_), .A3(new_n1712_), .ZN(new_n1713_));
  AND3_X1   g1521(.A1(new_n1700_), .A2(new_n1707_), .A3(new_n1642_), .ZN(new_n1714_));
  OAI211_X1 g1522(.A(new_n1505_), .B(new_n1511_), .C1(new_n1714_), .C2(new_n1708_), .ZN(new_n1715_));
  NAND2_X1  g1523(.A1(new_n1713_), .A2(new_n1715_), .ZN(new_n1716_));
  NOR2_X1   g1524(.A1(new_n648_), .A2(new_n616_), .ZN(new_n1717_));
  INV_X1    g1525(.A(new_n1717_), .ZN(new_n1718_));
  NAND3_X1  g1526(.A1(new_n1716_), .A2(KEYINPUT71), .A3(new_n1718_), .ZN(new_n1719_));
  NAND3_X1  g1527(.A1(new_n1713_), .A2(new_n1715_), .A3(new_n1717_), .ZN(new_n1720_));
  NAND3_X1  g1528(.A1(new_n1641_), .A2(new_n1719_), .A3(new_n1720_), .ZN(new_n1721_));
  AOI21_X1  g1529(.A(KEYINPUT71), .B1(new_n1716_), .B2(new_n1718_), .ZN(new_n1722_));
  OAI21_X1  g1530(.A(new_n1637_), .B1(new_n1721_), .B2(new_n1722_), .ZN(new_n1723_));
  NAND2_X1  g1531(.A1(new_n1716_), .A2(new_n1718_), .ZN(new_n1724_));
  NAND2_X1  g1532(.A1(new_n1724_), .A2(new_n1720_), .ZN(new_n1725_));
  NAND3_X1  g1533(.A1(new_n1725_), .A2(new_n1515_), .A3(new_n1524_), .ZN(new_n1726_));
  AND2_X1   g1534(.A1(new_n1713_), .A2(new_n1715_), .ZN(new_n1727_));
  AOI22_X1  g1535(.A1(new_n1524_), .A2(new_n1515_), .B1(new_n1727_), .B2(new_n1717_), .ZN(new_n1728_));
  INV_X1    g1536(.A(new_n1722_), .ZN(new_n1729_));
  NAND4_X1  g1537(.A1(new_n1728_), .A2(KEYINPUT72), .A3(new_n1729_), .A4(new_n1719_), .ZN(new_n1730_));
  NAND3_X1  g1538(.A1(new_n1723_), .A2(new_n1726_), .A3(new_n1730_), .ZN(new_n1731_));
  NOR2_X1   g1539(.A1(new_n539_), .A2(new_n774_), .ZN(new_n1732_));
  NAND2_X1  g1540(.A1(new_n1731_), .A2(new_n1732_), .ZN(new_n1733_));
  INV_X1    g1541(.A(KEYINPUT73), .ZN(new_n1734_));
  NAND2_X1  g1542(.A1(new_n1733_), .A2(new_n1734_), .ZN(new_n1735_));
  INV_X1    g1543(.A(new_n1732_), .ZN(new_n1736_));
  NAND4_X1  g1544(.A1(new_n1723_), .A2(new_n1730_), .A3(new_n1736_), .A4(new_n1726_), .ZN(new_n1737_));
  NAND2_X1  g1545(.A1(new_n1733_), .A2(new_n1737_), .ZN(new_n1738_));
  NAND3_X1  g1546(.A1(new_n1636_), .A2(new_n1735_), .A3(new_n1738_), .ZN(new_n1739_));
  NAND2_X1  g1547(.A1(new_n1536_), .A2(new_n1540_), .ZN(new_n1740_));
  AOI21_X1  g1548(.A(new_n1634_), .B1(new_n1740_), .B2(new_n1545_), .ZN(new_n1741_));
  OAI211_X1 g1549(.A(new_n1733_), .B(new_n1737_), .C1(new_n1741_), .C2(new_n1734_), .ZN(new_n1742_));
  NOR2_X1   g1550(.A1(new_n455_), .A2(new_n765_), .ZN(new_n1743_));
  INV_X1    g1551(.A(new_n1743_), .ZN(new_n1744_));
  AND3_X1   g1552(.A1(new_n1739_), .A2(new_n1742_), .A3(new_n1744_), .ZN(new_n1745_));
  AOI21_X1  g1553(.A(new_n1744_), .B1(new_n1739_), .B2(new_n1742_), .ZN(new_n1746_));
  OAI21_X1  g1554(.A(new_n1633_), .B1(new_n1745_), .B2(new_n1746_), .ZN(new_n1747_));
  NAND2_X1  g1555(.A1(new_n1739_), .A2(new_n1742_), .ZN(new_n1748_));
  NAND2_X1  g1556(.A1(new_n1748_), .A2(new_n1743_), .ZN(new_n1749_));
  NAND2_X1  g1557(.A1(new_n1562_), .A2(new_n1553_), .ZN(new_n1750_));
  NAND3_X1  g1558(.A1(new_n1739_), .A2(new_n1742_), .A3(new_n1744_), .ZN(new_n1751_));
  NAND3_X1  g1559(.A1(new_n1749_), .A2(new_n1750_), .A3(new_n1751_), .ZN(new_n1752_));
  NAND2_X1  g1560(.A1(G86gat), .A2(G460gat), .ZN(new_n1753_));
  NAND3_X1  g1561(.A1(new_n1747_), .A2(new_n1752_), .A3(new_n1753_), .ZN(new_n1754_));
  AOI21_X1  g1562(.A(new_n1753_), .B1(new_n1747_), .B2(new_n1752_), .ZN(new_n1755_));
  INV_X1    g1563(.A(new_n1755_), .ZN(new_n1756_));
  NAND3_X1  g1564(.A1(new_n1631_), .A2(new_n1754_), .A3(new_n1756_), .ZN(new_n1757_));
  AND3_X1   g1565(.A1(new_n1747_), .A2(new_n1752_), .A3(new_n1753_), .ZN(new_n1758_));
  OAI211_X1 g1566(.A(new_n1578_), .B(new_n1630_), .C1(new_n1758_), .C2(new_n1755_), .ZN(new_n1759_));
  NAND2_X1  g1567(.A1(new_n1757_), .A2(new_n1759_), .ZN(new_n1760_));
  NOR2_X1   g1568(.A1(new_n318_), .A2(new_n1215_), .ZN(new_n1761_));
  NAND2_X1  g1569(.A1(new_n1760_), .A2(new_n1761_), .ZN(new_n1762_));
  INV_X1    g1570(.A(new_n1761_), .ZN(new_n1763_));
  NAND3_X1  g1571(.A1(new_n1757_), .A2(new_n1759_), .A3(new_n1763_), .ZN(new_n1764_));
  AOI22_X1  g1572(.A1(new_n1582_), .A2(new_n1583_), .B1(G52gat), .B2(G477gat), .ZN(new_n1765_));
  NOR3_X1   g1573(.A1(new_n1568_), .A2(new_n1569_), .A3(new_n1574_), .ZN(new_n1766_));
  OAI211_X1 g1574(.A(new_n1762_), .B(new_n1764_), .C1(new_n1765_), .C2(new_n1766_), .ZN(new_n1767_));
  INV_X1    g1575(.A(new_n1766_), .ZN(new_n1768_));
  AND3_X1   g1576(.A1(new_n1757_), .A2(new_n1763_), .A3(new_n1759_), .ZN(new_n1769_));
  AOI21_X1  g1577(.A(new_n1763_), .B1(new_n1757_), .B2(new_n1759_), .ZN(new_n1770_));
  OAI211_X1 g1578(.A(new_n1580_), .B(new_n1768_), .C1(new_n1769_), .C2(new_n1770_), .ZN(new_n1771_));
  NAND2_X1  g1579(.A1(new_n1767_), .A2(new_n1771_), .ZN(new_n1772_));
  NOR2_X1   g1580(.A1(new_n214_), .A2(new_n1405_), .ZN(new_n1773_));
  NAND2_X1  g1581(.A1(new_n1772_), .A2(new_n1773_), .ZN(new_n1774_));
  INV_X1    g1582(.A(new_n1773_), .ZN(new_n1775_));
  NAND3_X1  g1583(.A1(new_n1767_), .A2(new_n1771_), .A3(new_n1775_), .ZN(new_n1776_));
  NAND2_X1  g1584(.A1(new_n1774_), .A2(new_n1776_), .ZN(new_n1777_));
  NAND3_X1  g1585(.A1(new_n1767_), .A2(new_n1771_), .A3(new_n1773_), .ZN(new_n1778_));
  INV_X1    g1586(.A(KEYINPUT74), .ZN(new_n1779_));
  AND2_X1   g1587(.A1(new_n1778_), .A2(new_n1779_), .ZN(new_n1780_));
  AOI21_X1  g1588(.A(new_n1596_), .B1(new_n1402_), .B2(new_n1586_), .ZN(new_n1781_));
  AOI21_X1  g1589(.A(new_n1781_), .B1(new_n1609_), .B2(new_n1610_), .ZN(new_n1782_));
  OAI21_X1  g1590(.A(new_n1777_), .B1(new_n1780_), .B2(new_n1782_), .ZN(new_n1783_));
  INV_X1    g1591(.A(new_n1781_), .ZN(new_n1784_));
  OAI21_X1  g1592(.A(new_n1784_), .B1(new_n1598_), .B2(new_n1599_), .ZN(new_n1785_));
  NAND2_X1  g1593(.A1(new_n1778_), .A2(new_n1779_), .ZN(new_n1786_));
  NAND4_X1  g1594(.A1(new_n1785_), .A2(new_n1786_), .A3(new_n1776_), .A4(new_n1774_), .ZN(new_n1787_));
  NAND2_X1  g1595(.A1(new_n1783_), .A2(new_n1787_), .ZN(new_n1788_));
  NOR2_X1   g1596(.A1(new_n213_), .A2(new_n1417_), .ZN(new_n1789_));
  NAND2_X1  g1597(.A1(new_n1788_), .A2(new_n1789_), .ZN(new_n1790_));
  NAND2_X1  g1598(.A1(G35gat), .A2(G511gat), .ZN(new_n1791_));
  NAND3_X1  g1599(.A1(new_n1783_), .A2(new_n1787_), .A3(new_n1791_), .ZN(new_n1792_));
  AND3_X1   g1600(.A1(new_n1629_), .A2(new_n1790_), .A3(new_n1792_), .ZN(new_n1793_));
  AOI21_X1  g1601(.A(new_n1629_), .B1(new_n1790_), .B2(new_n1792_), .ZN(new_n1794_));
  NOR2_X1   g1602(.A1(new_n196_), .A2(new_n1622_), .ZN(new_n1795_));
  NOR3_X1   g1603(.A1(new_n1793_), .A2(new_n1794_), .A3(new_n1795_), .ZN(new_n1796_));
  INV_X1    g1604(.A(new_n1795_), .ZN(new_n1797_));
  NAND2_X1  g1605(.A1(new_n1790_), .A2(new_n1792_), .ZN(new_n1798_));
  AND2_X1   g1606(.A1(new_n1616_), .A2(new_n1628_), .ZN(new_n1799_));
  NAND2_X1  g1607(.A1(new_n1798_), .A2(new_n1799_), .ZN(new_n1800_));
  NAND3_X1  g1608(.A1(new_n1629_), .A2(new_n1790_), .A3(new_n1792_), .ZN(new_n1801_));
  AOI21_X1  g1609(.A(new_n1797_), .B1(new_n1800_), .B2(new_n1801_), .ZN(new_n1802_));
  NOR2_X1   g1610(.A1(new_n1796_), .A2(new_n1802_), .ZN(new_n1803_));
  INV_X1    g1611(.A(new_n1623_), .ZN(new_n1804_));
  AOI21_X1  g1612(.A(new_n1618_), .B1(new_n1804_), .B2(new_n1620_), .ZN(new_n1805_));
  XNOR2_X1  g1613(.A(new_n1803_), .B(new_n1805_), .ZN(G6150gat));
  AOI21_X1  g1614(.A(new_n1793_), .B1(new_n1797_), .B2(new_n1800_), .ZN(new_n1807_));
  NAND3_X1  g1615(.A1(new_n1785_), .A2(new_n1776_), .A3(new_n1774_), .ZN(new_n1808_));
  NAND2_X1  g1616(.A1(new_n1776_), .A2(KEYINPUT75), .ZN(new_n1809_));
  NOR2_X1   g1617(.A1(new_n312_), .A2(new_n1215_), .ZN(new_n1810_));
  NOR2_X1   g1618(.A1(new_n539_), .A2(new_n765_), .ZN(new_n1811_));
  INV_X1    g1619(.A(new_n1811_), .ZN(new_n1812_));
  NAND2_X1  g1620(.A1(new_n1727_), .A2(new_n1718_), .ZN(new_n1813_));
  INV_X1    g1621(.A(KEYINPUT78), .ZN(new_n1814_));
  AOI211_X1 g1622(.A(new_n1708_), .B(new_n1714_), .C1(new_n1711_), .C2(new_n1814_), .ZN(new_n1815_));
  OAI21_X1  g1623(.A(new_n1815_), .B1(new_n1814_), .B2(new_n1711_), .ZN(new_n1816_));
  NAND2_X1  g1624(.A1(new_n1813_), .A2(new_n1816_), .ZN(new_n1817_));
  NAND2_X1  g1625(.A1(new_n1712_), .A2(new_n1707_), .ZN(new_n1818_));
  INV_X1    g1626(.A(new_n1818_), .ZN(new_n1819_));
  INV_X1    g1627(.A(KEYINPUT79), .ZN(new_n1820_));
  AOI22_X1  g1628(.A1(new_n1653_), .A2(new_n1672_), .B1(new_n1649_), .B2(new_n1675_), .ZN(new_n1821_));
  NAND2_X1  g1629(.A1(new_n1671_), .A2(new_n1669_), .ZN(new_n1822_));
  INV_X1    g1630(.A(G256gat), .ZN(new_n1823_));
  NAND2_X1  g1631(.A1(new_n1262_), .A2(G273gat), .ZN(new_n1824_));
  AOI21_X1  g1632(.A(new_n1823_), .B1(new_n1824_), .B2(new_n245_), .ZN(new_n1825_));
  NAND2_X1  g1633(.A1(new_n1658_), .A2(G290gat), .ZN(new_n1826_));
  NAND2_X1  g1634(.A1(new_n1825_), .A2(new_n1826_), .ZN(new_n1827_));
  NAND2_X1  g1635(.A1(G239gat), .A2(G324gat), .ZN(new_n1828_));
  XNOR2_X1  g1636(.A(new_n1827_), .B(new_n1828_), .ZN(new_n1829_));
  INV_X1    g1637(.A(new_n1829_), .ZN(new_n1830_));
  NOR2_X1   g1638(.A1(new_n1822_), .A2(new_n1830_), .ZN(new_n1831_));
  OAI21_X1  g1639(.A(new_n1671_), .B1(new_n1665_), .B2(new_n1666_), .ZN(new_n1832_));
  AOI21_X1  g1640(.A(new_n1831_), .B1(new_n1832_), .B2(new_n1830_), .ZN(new_n1833_));
  NOR2_X1   g1641(.A1(new_n1437_), .A2(new_n261_), .ZN(new_n1834_));
  NOR2_X1   g1642(.A1(new_n1822_), .A2(new_n1829_), .ZN(new_n1835_));
  NOR2_X1   g1643(.A1(new_n1835_), .A2(new_n1834_), .ZN(new_n1836_));
  NAND2_X1  g1644(.A1(new_n1832_), .A2(new_n1829_), .ZN(new_n1837_));
  AOI22_X1  g1645(.A1(new_n1833_), .A2(new_n1834_), .B1(new_n1836_), .B2(new_n1837_), .ZN(new_n1838_));
  INV_X1    g1646(.A(new_n1838_), .ZN(new_n1839_));
  OR2_X1    g1647(.A1(new_n1821_), .A2(new_n1839_), .ZN(new_n1840_));
  NOR2_X1   g1648(.A1(new_n302_), .A2(new_n942_), .ZN(new_n1841_));
  INV_X1    g1649(.A(new_n1841_), .ZN(new_n1842_));
  NAND2_X1  g1650(.A1(new_n1821_), .A2(new_n1839_), .ZN(new_n1843_));
  NAND3_X1  g1651(.A1(new_n1840_), .A2(new_n1842_), .A3(new_n1843_), .ZN(new_n1844_));
  AOI221_X4 g1652(.A(new_n1838_), .B1(new_n1649_), .B2(new_n1675_), .C1(new_n1653_), .C2(new_n1672_), .ZN(new_n1845_));
  NOR2_X1   g1653(.A1(new_n1821_), .A2(new_n1839_), .ZN(new_n1846_));
  OAI21_X1  g1654(.A(new_n1841_), .B1(new_n1845_), .B2(new_n1846_), .ZN(new_n1847_));
  NAND2_X1  g1655(.A1(new_n1844_), .A2(new_n1847_), .ZN(new_n1848_));
  NAND3_X1  g1656(.A1(new_n1848_), .A2(new_n1687_), .A3(new_n1694_), .ZN(new_n1849_));
  AOI21_X1  g1657(.A(new_n1685_), .B1(new_n1683_), .B2(new_n1686_), .ZN(new_n1850_));
  OAI21_X1  g1658(.A(new_n1687_), .B1(new_n1850_), .B2(new_n1681_), .ZN(new_n1851_));
  NAND3_X1  g1659(.A1(new_n1851_), .A2(new_n1844_), .A3(new_n1847_), .ZN(new_n1852_));
  NOR2_X1   g1660(.A1(new_n1092_), .A2(new_n356_), .ZN(new_n1853_));
  INV_X1    g1661(.A(new_n1853_), .ZN(new_n1854_));
  AND3_X1   g1662(.A1(new_n1849_), .A2(new_n1852_), .A3(new_n1854_), .ZN(new_n1855_));
  AOI21_X1  g1663(.A(new_n1854_), .B1(new_n1849_), .B2(new_n1852_), .ZN(new_n1856_));
  OAI21_X1  g1664(.A(new_n1820_), .B1(new_n1855_), .B2(new_n1856_), .ZN(new_n1857_));
  NAND2_X1  g1665(.A1(new_n1706_), .A2(new_n1695_), .ZN(new_n1858_));
  NAND3_X1  g1666(.A1(new_n1849_), .A2(new_n1852_), .A3(KEYINPUT79), .ZN(new_n1859_));
  NAND3_X1  g1667(.A1(new_n1857_), .A2(new_n1858_), .A3(new_n1859_), .ZN(new_n1860_));
  NOR2_X1   g1668(.A1(new_n946_), .A2(new_n867_), .ZN(new_n1861_));
  INV_X1    g1669(.A(new_n1861_), .ZN(new_n1862_));
  OAI211_X1 g1670(.A(new_n1695_), .B(new_n1706_), .C1(new_n1855_), .C2(new_n1856_), .ZN(new_n1863_));
  NAND3_X1  g1671(.A1(new_n1860_), .A2(new_n1862_), .A3(new_n1863_), .ZN(new_n1864_));
  INV_X1    g1672(.A(new_n1864_), .ZN(new_n1865_));
  AOI21_X1  g1673(.A(new_n1862_), .B1(new_n1860_), .B2(new_n1863_), .ZN(new_n1866_));
  OAI21_X1  g1674(.A(new_n1819_), .B1(new_n1865_), .B2(new_n1866_), .ZN(new_n1867_));
  NOR2_X1   g1675(.A1(new_n957_), .A2(new_n616_), .ZN(new_n1868_));
  NAND2_X1  g1676(.A1(new_n1860_), .A2(new_n1863_), .ZN(new_n1869_));
  NAND2_X1  g1677(.A1(new_n1869_), .A2(new_n1861_), .ZN(new_n1870_));
  NAND3_X1  g1678(.A1(new_n1870_), .A2(new_n1818_), .A3(new_n1864_), .ZN(new_n1871_));
  NAND3_X1  g1679(.A1(new_n1867_), .A2(new_n1868_), .A3(new_n1871_), .ZN(new_n1872_));
  AOI21_X1  g1680(.A(new_n1868_), .B1(new_n1867_), .B2(new_n1871_), .ZN(new_n1873_));
  OAI21_X1  g1681(.A(new_n1872_), .B1(new_n1873_), .B2(KEYINPUT80), .ZN(new_n1874_));
  INV_X1    g1682(.A(KEYINPUT80), .ZN(new_n1875_));
  AOI211_X1 g1683(.A(new_n1875_), .B(new_n1868_), .C1(new_n1867_), .C2(new_n1871_), .ZN(new_n1876_));
  OAI21_X1  g1684(.A(new_n1817_), .B1(new_n1874_), .B2(new_n1876_), .ZN(new_n1877_));
  INV_X1    g1685(.A(new_n1873_), .ZN(new_n1878_));
  NAND4_X1  g1686(.A1(new_n1878_), .A2(new_n1813_), .A3(new_n1816_), .A4(new_n1872_), .ZN(new_n1879_));
  NAND2_X1  g1687(.A1(new_n1877_), .A2(new_n1879_), .ZN(new_n1880_));
  NOR2_X1   g1688(.A1(new_n648_), .A2(new_n774_), .ZN(new_n1881_));
  INV_X1    g1689(.A(new_n1881_), .ZN(new_n1882_));
  NAND2_X1  g1690(.A1(new_n1880_), .A2(new_n1882_), .ZN(new_n1883_));
  NAND3_X1  g1691(.A1(new_n1877_), .A2(new_n1881_), .A3(new_n1879_), .ZN(new_n1884_));
  NAND2_X1  g1692(.A1(new_n1883_), .A2(new_n1884_), .ZN(new_n1885_));
  AND2_X1   g1693(.A1(new_n1725_), .A2(new_n1641_), .ZN(new_n1886_));
  NAND2_X1  g1694(.A1(new_n1731_), .A2(new_n1736_), .ZN(new_n1887_));
  AOI21_X1  g1695(.A(new_n1886_), .B1(new_n1887_), .B2(KEYINPUT82), .ZN(new_n1888_));
  INV_X1    g1696(.A(KEYINPUT82), .ZN(new_n1889_));
  NAND3_X1  g1697(.A1(new_n1731_), .A2(new_n1889_), .A3(new_n1736_), .ZN(new_n1890_));
  AOI21_X1  g1698(.A(new_n1885_), .B1(new_n1888_), .B2(new_n1890_), .ZN(new_n1891_));
  INV_X1    g1699(.A(KEYINPUT81), .ZN(new_n1892_));
  NAND3_X1  g1700(.A1(new_n1883_), .A2(new_n1892_), .A3(new_n1884_), .ZN(new_n1893_));
  NAND3_X1  g1701(.A1(new_n1880_), .A2(KEYINPUT81), .A3(new_n1882_), .ZN(new_n1894_));
  AOI21_X1  g1702(.A(new_n1886_), .B1(new_n1731_), .B2(new_n1736_), .ZN(new_n1895_));
  AND3_X1   g1703(.A1(new_n1893_), .A2(new_n1894_), .A3(new_n1895_), .ZN(new_n1896_));
  OAI21_X1  g1704(.A(new_n1812_), .B1(new_n1891_), .B2(new_n1896_), .ZN(new_n1897_));
  NAND3_X1  g1705(.A1(new_n1893_), .A2(new_n1894_), .A3(new_n1895_), .ZN(new_n1898_));
  AND3_X1   g1706(.A1(new_n1731_), .A2(new_n1889_), .A3(new_n1736_), .ZN(new_n1899_));
  AOI21_X1  g1707(.A(new_n1889_), .B1(new_n1731_), .B2(new_n1736_), .ZN(new_n1900_));
  NOR3_X1   g1708(.A1(new_n1899_), .A2(new_n1900_), .A3(new_n1886_), .ZN(new_n1901_));
  OAI211_X1 g1709(.A(new_n1811_), .B(new_n1898_), .C1(new_n1901_), .C2(new_n1885_), .ZN(new_n1902_));
  NAND2_X1  g1710(.A1(new_n1738_), .A2(KEYINPUT77), .ZN(new_n1903_));
  INV_X1    g1711(.A(KEYINPUT77), .ZN(new_n1904_));
  NAND3_X1  g1712(.A1(new_n1733_), .A2(new_n1904_), .A3(new_n1737_), .ZN(new_n1905_));
  NAND3_X1  g1713(.A1(new_n1903_), .A2(new_n1636_), .A3(new_n1905_), .ZN(new_n1906_));
  NAND2_X1  g1714(.A1(new_n1906_), .A2(KEYINPUT76), .ZN(new_n1907_));
  NAND3_X1  g1715(.A1(new_n1897_), .A2(new_n1902_), .A3(new_n1907_), .ZN(new_n1908_));
  NAND2_X1  g1716(.A1(new_n1751_), .A2(new_n1906_), .ZN(new_n1909_));
  INV_X1    g1717(.A(new_n1909_), .ZN(new_n1910_));
  NAND2_X1  g1718(.A1(new_n1908_), .A2(new_n1910_), .ZN(new_n1911_));
  NOR2_X1   g1719(.A1(new_n455_), .A2(new_n1055_), .ZN(new_n1912_));
  INV_X1    g1720(.A(new_n1912_), .ZN(new_n1913_));
  NAND4_X1  g1721(.A1(new_n1909_), .A2(new_n1897_), .A3(new_n1902_), .A4(new_n1907_), .ZN(new_n1914_));
  AND3_X1   g1722(.A1(new_n1911_), .A2(new_n1913_), .A3(new_n1914_), .ZN(new_n1915_));
  AOI21_X1  g1723(.A(new_n1913_), .B1(new_n1911_), .B2(new_n1914_), .ZN(new_n1916_));
  NOR3_X1   g1724(.A1(new_n1745_), .A2(new_n1633_), .A3(new_n1746_), .ZN(new_n1917_));
  AOI21_X1  g1725(.A(new_n1917_), .B1(new_n1753_), .B2(new_n1747_), .ZN(new_n1918_));
  NOR3_X1   g1726(.A1(new_n1915_), .A2(new_n1916_), .A3(new_n1918_), .ZN(new_n1919_));
  NAND2_X1  g1727(.A1(new_n1754_), .A2(new_n1752_), .ZN(new_n1920_));
  NAND2_X1  g1728(.A1(new_n1911_), .A2(new_n1914_), .ZN(new_n1921_));
  NAND2_X1  g1729(.A1(new_n1921_), .A2(new_n1912_), .ZN(new_n1922_));
  NAND3_X1  g1730(.A1(new_n1911_), .A2(new_n1913_), .A3(new_n1914_), .ZN(new_n1923_));
  AOI21_X1  g1731(.A(new_n1920_), .B1(new_n1922_), .B2(new_n1923_), .ZN(new_n1924_));
  OAI21_X1  g1732(.A(new_n1810_), .B1(new_n1919_), .B2(new_n1924_), .ZN(new_n1925_));
  OAI21_X1  g1733(.A(new_n1918_), .B1(new_n1915_), .B2(new_n1916_), .ZN(new_n1926_));
  NAND3_X1  g1734(.A1(new_n1922_), .A2(new_n1920_), .A3(new_n1923_), .ZN(new_n1927_));
  INV_X1    g1735(.A(new_n1810_), .ZN(new_n1928_));
  NAND3_X1  g1736(.A1(new_n1926_), .A2(new_n1927_), .A3(new_n1928_), .ZN(new_n1929_));
  NAND2_X1  g1737(.A1(new_n1925_), .A2(new_n1929_), .ZN(new_n1930_));
  NAND3_X1  g1738(.A1(new_n1930_), .A2(new_n1757_), .A3(new_n1764_), .ZN(new_n1931_));
  NOR2_X1   g1739(.A1(new_n318_), .A2(new_n1405_), .ZN(new_n1932_));
  INV_X1    g1740(.A(new_n1932_), .ZN(new_n1933_));
  NAND2_X1  g1741(.A1(new_n1764_), .A2(new_n1757_), .ZN(new_n1934_));
  NAND3_X1  g1742(.A1(new_n1925_), .A2(new_n1934_), .A3(new_n1929_), .ZN(new_n1935_));
  NAND3_X1  g1743(.A1(new_n1931_), .A2(new_n1933_), .A3(new_n1935_), .ZN(new_n1936_));
  AND3_X1   g1744(.A1(new_n1925_), .A2(new_n1934_), .A3(new_n1929_), .ZN(new_n1937_));
  AOI21_X1  g1745(.A(new_n1934_), .B1(new_n1925_), .B2(new_n1929_), .ZN(new_n1938_));
  OAI21_X1  g1746(.A(new_n1932_), .B1(new_n1937_), .B2(new_n1938_), .ZN(new_n1939_));
  NAND3_X1  g1747(.A1(new_n1809_), .A2(new_n1936_), .A3(new_n1939_), .ZN(new_n1940_));
  NAND2_X1  g1748(.A1(new_n1776_), .A2(new_n1767_), .ZN(new_n1941_));
  INV_X1    g1749(.A(new_n1941_), .ZN(new_n1942_));
  NAND2_X1  g1750(.A1(new_n1940_), .A2(new_n1942_), .ZN(new_n1943_));
  NOR2_X1   g1751(.A1(new_n214_), .A2(new_n1417_), .ZN(new_n1944_));
  INV_X1    g1752(.A(new_n1944_), .ZN(new_n1945_));
  NAND4_X1  g1753(.A1(new_n1941_), .A2(new_n1809_), .A3(new_n1936_), .A4(new_n1939_), .ZN(new_n1946_));
  AND3_X1   g1754(.A1(new_n1943_), .A2(new_n1945_), .A3(new_n1946_), .ZN(new_n1947_));
  AOI21_X1  g1755(.A(new_n1945_), .B1(new_n1943_), .B2(new_n1946_), .ZN(new_n1948_));
  OAI211_X1 g1756(.A(new_n1792_), .B(new_n1808_), .C1(new_n1947_), .C2(new_n1948_), .ZN(new_n1949_));
  NAND2_X1  g1757(.A1(new_n1792_), .A2(new_n1808_), .ZN(new_n1950_));
  NAND2_X1  g1758(.A1(new_n1943_), .A2(new_n1946_), .ZN(new_n1951_));
  NAND2_X1  g1759(.A1(new_n1951_), .A2(new_n1944_), .ZN(new_n1952_));
  NAND3_X1  g1760(.A1(new_n1943_), .A2(new_n1945_), .A3(new_n1946_), .ZN(new_n1953_));
  NAND3_X1  g1761(.A1(new_n1950_), .A2(new_n1952_), .A3(new_n1953_), .ZN(new_n1954_));
  NOR2_X1   g1762(.A1(new_n213_), .A2(new_n1622_), .ZN(new_n1955_));
  XNOR2_X1  g1763(.A(new_n1955_), .B(KEYINPUT83), .ZN(new_n1956_));
  INV_X1    g1764(.A(new_n1956_), .ZN(new_n1957_));
  AND3_X1   g1765(.A1(new_n1949_), .A2(new_n1954_), .A3(new_n1957_), .ZN(new_n1958_));
  AOI21_X1  g1766(.A(new_n1957_), .B1(new_n1949_), .B2(new_n1954_), .ZN(new_n1959_));
  OAI21_X1  g1767(.A(new_n1807_), .B1(new_n1958_), .B2(new_n1959_), .ZN(new_n1960_));
  NAND2_X1  g1768(.A1(new_n1949_), .A2(new_n1954_), .ZN(new_n1961_));
  NAND2_X1  g1769(.A1(new_n1961_), .A2(new_n1956_), .ZN(new_n1962_));
  OAI21_X1  g1770(.A(new_n1801_), .B1(new_n1794_), .B2(new_n1795_), .ZN(new_n1963_));
  NAND3_X1  g1771(.A1(new_n1949_), .A2(new_n1954_), .A3(new_n1955_), .ZN(new_n1964_));
  NAND3_X1  g1772(.A1(new_n1962_), .A2(new_n1963_), .A3(new_n1964_), .ZN(new_n1965_));
  NAND2_X1  g1773(.A1(new_n1960_), .A2(new_n1965_), .ZN(new_n1966_));
  OAI21_X1  g1774(.A(new_n1805_), .B1(new_n1796_), .B2(new_n1802_), .ZN(new_n1967_));
  XNOR2_X1  g1775(.A(new_n1966_), .B(new_n1967_), .ZN(G6160gat));
  NAND3_X1  g1776(.A1(new_n1949_), .A2(new_n1954_), .A3(new_n1957_), .ZN(new_n1969_));
  AOI21_X1  g1777(.A(new_n1807_), .B1(new_n1962_), .B2(new_n1969_), .ZN(new_n1970_));
  AOI21_X1  g1778(.A(new_n1970_), .B1(new_n1966_), .B2(new_n1967_), .ZN(new_n1971_));
  AOI21_X1  g1779(.A(new_n1950_), .B1(new_n1953_), .B2(new_n1952_), .ZN(new_n1972_));
  OAI21_X1  g1780(.A(new_n1954_), .B1(new_n1972_), .B2(new_n1955_), .ZN(new_n1973_));
  INV_X1    g1781(.A(KEYINPUT88), .ZN(new_n1974_));
  AOI21_X1  g1782(.A(new_n1937_), .B1(new_n1931_), .B2(new_n1933_), .ZN(new_n1975_));
  AOI21_X1  g1783(.A(new_n1919_), .B1(new_n1928_), .B2(new_n1926_), .ZN(new_n1976_));
  NAND3_X1  g1784(.A1(new_n1909_), .A2(new_n1897_), .A3(new_n1902_), .ZN(new_n1977_));
  AND2_X1   g1785(.A1(new_n1923_), .A2(new_n1977_), .ZN(new_n1978_));
  INV_X1    g1786(.A(KEYINPUT87), .ZN(new_n1979_));
  NAND2_X1  g1787(.A1(new_n1977_), .A2(new_n1979_), .ZN(new_n1980_));
  AND2_X1   g1788(.A1(new_n1893_), .A2(new_n1894_), .ZN(new_n1981_));
  NAND2_X1  g1789(.A1(new_n1887_), .A2(KEYINPUT82), .ZN(new_n1982_));
  INV_X1    g1790(.A(new_n1886_), .ZN(new_n1983_));
  NAND3_X1  g1791(.A1(new_n1982_), .A2(new_n1890_), .A3(new_n1983_), .ZN(new_n1984_));
  NAND2_X1  g1792(.A1(new_n1981_), .A2(new_n1984_), .ZN(new_n1985_));
  NOR2_X1   g1793(.A1(new_n648_), .A2(new_n765_), .ZN(new_n1986_));
  NOR2_X1   g1794(.A1(new_n946_), .A2(new_n616_), .ZN(new_n1987_));
  NOR2_X1   g1795(.A1(new_n1092_), .A2(new_n867_), .ZN(new_n1988_));
  INV_X1    g1796(.A(KEYINPUT85), .ZN(new_n1989_));
  NAND2_X1  g1797(.A1(new_n1988_), .A2(new_n1989_), .ZN(new_n1990_));
  INV_X1    g1798(.A(new_n1988_), .ZN(new_n1991_));
  NAND2_X1  g1799(.A1(new_n1991_), .A2(KEYINPUT85), .ZN(new_n1992_));
  INV_X1    g1800(.A(new_n1837_), .ZN(new_n1993_));
  NOR2_X1   g1801(.A1(new_n1993_), .A2(new_n1836_), .ZN(new_n1994_));
  INV_X1    g1802(.A(new_n1828_), .ZN(new_n1995_));
  OAI21_X1  g1803(.A(new_n1825_), .B1(new_n1827_), .B2(new_n1995_), .ZN(new_n1996_));
  OR2_X1    g1804(.A1(new_n1996_), .A2(new_n232_), .ZN(new_n1997_));
  OAI21_X1  g1805(.A(new_n1996_), .B1(new_n1823_), .B2(new_n232_), .ZN(new_n1998_));
  NAND2_X1  g1806(.A1(new_n1997_), .A2(new_n1998_), .ZN(new_n1999_));
  NAND2_X1  g1807(.A1(G239gat), .A2(G341gat), .ZN(new_n2000_));
  XOR2_X1   g1808(.A(new_n1999_), .B(new_n2000_), .Z(new_n2001_));
  NAND2_X1  g1809(.A1(new_n1994_), .A2(new_n2001_), .ZN(new_n2002_));
  NAND2_X1  g1810(.A1(new_n1832_), .A2(new_n1830_), .ZN(new_n2003_));
  OAI21_X1  g1811(.A(new_n2003_), .B1(new_n1830_), .B2(new_n1822_), .ZN(new_n2004_));
  INV_X1    g1812(.A(new_n1834_), .ZN(new_n2005_));
  AOI21_X1  g1813(.A(new_n1993_), .B1(new_n2004_), .B2(new_n2005_), .ZN(new_n2006_));
  OAI21_X1  g1814(.A(new_n2002_), .B1(new_n2006_), .B2(new_n2001_), .ZN(new_n2007_));
  NAND2_X1  g1815(.A1(new_n348_), .A2(G222gat), .ZN(new_n2008_));
  XOR2_X1   g1816(.A(new_n2007_), .B(new_n2008_), .Z(new_n2009_));
  AOI21_X1  g1817(.A(new_n1846_), .B1(new_n1842_), .B2(new_n1843_), .ZN(new_n2010_));
  XNOR2_X1  g1818(.A(new_n2009_), .B(new_n2010_), .ZN(new_n2011_));
  NOR2_X1   g1819(.A1(new_n942_), .A2(new_n356_), .ZN(new_n2012_));
  XOR2_X1   g1820(.A(new_n2011_), .B(new_n2012_), .Z(new_n2013_));
  INV_X1    g1821(.A(KEYINPUT84), .ZN(new_n2014_));
  NAND2_X1  g1822(.A1(new_n1849_), .A2(new_n1852_), .ZN(new_n2015_));
  OAI211_X1 g1823(.A(new_n2014_), .B(new_n1852_), .C1(new_n2015_), .C2(new_n1853_), .ZN(new_n2016_));
  OAI21_X1  g1824(.A(new_n1852_), .B1(new_n2015_), .B2(new_n1853_), .ZN(new_n2017_));
  NAND2_X1  g1825(.A1(new_n2017_), .A2(KEYINPUT84), .ZN(new_n2018_));
  AOI21_X1  g1826(.A(new_n2013_), .B1(new_n2016_), .B2(new_n2018_), .ZN(new_n2019_));
  XNOR2_X1  g1827(.A(new_n2011_), .B(new_n2012_), .ZN(new_n2020_));
  AOI21_X1  g1828(.A(new_n2020_), .B1(KEYINPUT84), .B2(new_n2017_), .ZN(new_n2021_));
  OAI211_X1 g1829(.A(new_n1990_), .B(new_n1992_), .C1(new_n2019_), .C2(new_n2021_), .ZN(new_n2022_));
  NAND2_X1  g1830(.A1(new_n2018_), .A2(new_n2016_), .ZN(new_n2023_));
  NAND2_X1  g1831(.A1(new_n2023_), .A2(new_n2020_), .ZN(new_n2024_));
  NAND2_X1  g1832(.A1(new_n2013_), .A2(new_n2018_), .ZN(new_n2025_));
  NAND4_X1  g1833(.A1(new_n2024_), .A2(new_n1989_), .A3(new_n1988_), .A4(new_n2025_), .ZN(new_n2026_));
  NAND2_X1  g1834(.A1(new_n1864_), .A2(new_n1860_), .ZN(new_n2027_));
  AND3_X1   g1835(.A1(new_n2022_), .A2(new_n2026_), .A3(new_n2027_), .ZN(new_n2028_));
  AOI21_X1  g1836(.A(new_n2027_), .B1(new_n2022_), .B2(new_n2026_), .ZN(new_n2029_));
  OAI21_X1  g1837(.A(new_n1987_), .B1(new_n2028_), .B2(new_n2029_), .ZN(new_n2030_));
  NAND2_X1  g1838(.A1(new_n2022_), .A2(new_n2026_), .ZN(new_n2031_));
  INV_X1    g1839(.A(new_n2027_), .ZN(new_n2032_));
  NAND2_X1  g1840(.A1(new_n2031_), .A2(new_n2032_), .ZN(new_n2033_));
  INV_X1    g1841(.A(new_n1987_), .ZN(new_n2034_));
  NAND3_X1  g1842(.A1(new_n2022_), .A2(new_n2026_), .A3(new_n2027_), .ZN(new_n2035_));
  NAND3_X1  g1843(.A1(new_n2033_), .A2(new_n2034_), .A3(new_n2035_), .ZN(new_n2036_));
  NAND2_X1  g1844(.A1(new_n2030_), .A2(new_n2036_), .ZN(new_n2037_));
  OAI211_X1 g1845(.A(new_n1867_), .B(new_n1871_), .C1(new_n957_), .C2(new_n616_), .ZN(new_n2038_));
  XNOR2_X1  g1846(.A(new_n1871_), .B(KEYINPUT86), .ZN(new_n2039_));
  NAND3_X1  g1847(.A1(new_n2037_), .A2(new_n2038_), .A3(new_n2039_), .ZN(new_n2040_));
  NAND2_X1  g1848(.A1(new_n2039_), .A2(new_n2038_), .ZN(new_n2041_));
  NAND3_X1  g1849(.A1(new_n2041_), .A2(new_n2036_), .A3(new_n2030_), .ZN(new_n2042_));
  NAND2_X1  g1850(.A1(new_n2040_), .A2(new_n2042_), .ZN(new_n2043_));
  NOR2_X1   g1851(.A1(new_n957_), .A2(new_n774_), .ZN(new_n2044_));
  NAND2_X1  g1852(.A1(new_n2043_), .A2(new_n2044_), .ZN(new_n2045_));
  OAI211_X1 g1853(.A(new_n2040_), .B(new_n2042_), .C1(new_n957_), .C2(new_n774_), .ZN(new_n2046_));
  NOR2_X1   g1854(.A1(new_n1817_), .A2(new_n1873_), .ZN(new_n2047_));
  AOI22_X1  g1855(.A1(new_n1877_), .A2(new_n1881_), .B1(new_n2047_), .B2(new_n1872_), .ZN(new_n2048_));
  AND3_X1   g1856(.A1(new_n2045_), .A2(new_n2046_), .A3(new_n2048_), .ZN(new_n2049_));
  AOI21_X1  g1857(.A(new_n2048_), .B1(new_n2045_), .B2(new_n2046_), .ZN(new_n2050_));
  OAI21_X1  g1858(.A(new_n1986_), .B1(new_n2049_), .B2(new_n2050_), .ZN(new_n2051_));
  NAND2_X1  g1859(.A1(new_n2045_), .A2(new_n2046_), .ZN(new_n2052_));
  INV_X1    g1860(.A(new_n2048_), .ZN(new_n2053_));
  NAND2_X1  g1861(.A1(new_n2052_), .A2(new_n2053_), .ZN(new_n2054_));
  INV_X1    g1862(.A(new_n1986_), .ZN(new_n2055_));
  NAND3_X1  g1863(.A1(new_n2045_), .A2(new_n2046_), .A3(new_n2048_), .ZN(new_n2056_));
  NAND3_X1  g1864(.A1(new_n2054_), .A2(new_n2055_), .A3(new_n2056_), .ZN(new_n2057_));
  NAND2_X1  g1865(.A1(new_n2051_), .A2(new_n2057_), .ZN(new_n2058_));
  AND3_X1   g1866(.A1(new_n1897_), .A2(new_n1985_), .A3(new_n2058_), .ZN(new_n2059_));
  AOI21_X1  g1867(.A(new_n2058_), .B1(new_n1897_), .B2(new_n1985_), .ZN(new_n2060_));
  NOR2_X1   g1868(.A1(new_n539_), .A2(new_n1055_), .ZN(new_n2061_));
  NOR3_X1   g1869(.A1(new_n2059_), .A2(new_n2060_), .A3(new_n2061_), .ZN(new_n2062_));
  INV_X1    g1870(.A(new_n2061_), .ZN(new_n2063_));
  INV_X1    g1871(.A(new_n2058_), .ZN(new_n2064_));
  INV_X1    g1872(.A(new_n1885_), .ZN(new_n2065_));
  NAND2_X1  g1873(.A1(new_n1984_), .A2(new_n2065_), .ZN(new_n2066_));
  AOI21_X1  g1874(.A(new_n1811_), .B1(new_n2066_), .B2(new_n1898_), .ZN(new_n2067_));
  INV_X1    g1875(.A(new_n1985_), .ZN(new_n2068_));
  OAI21_X1  g1876(.A(new_n2064_), .B1(new_n2067_), .B2(new_n2068_), .ZN(new_n2069_));
  NAND3_X1  g1877(.A1(new_n1897_), .A2(new_n1985_), .A3(new_n2058_), .ZN(new_n2070_));
  AOI21_X1  g1878(.A(new_n2063_), .B1(new_n2069_), .B2(new_n2070_), .ZN(new_n2071_));
  OAI21_X1  g1879(.A(new_n1980_), .B1(new_n2062_), .B2(new_n2071_), .ZN(new_n2072_));
  NAND2_X1  g1880(.A1(new_n1978_), .A2(new_n2072_), .ZN(new_n2073_));
  NOR2_X1   g1881(.A1(new_n455_), .A2(new_n1215_), .ZN(new_n2074_));
  NAND2_X1  g1882(.A1(new_n1923_), .A2(new_n1977_), .ZN(new_n2075_));
  OAI21_X1  g1883(.A(new_n2061_), .B1(new_n2059_), .B2(new_n2060_), .ZN(new_n2076_));
  NAND3_X1  g1884(.A1(new_n2069_), .A2(new_n2063_), .A3(new_n2070_), .ZN(new_n2077_));
  NAND2_X1  g1885(.A1(new_n2076_), .A2(new_n2077_), .ZN(new_n2078_));
  NAND3_X1  g1886(.A1(new_n2075_), .A2(new_n2078_), .A3(new_n1980_), .ZN(new_n2079_));
  AND3_X1   g1887(.A1(new_n2073_), .A2(new_n2074_), .A3(new_n2079_), .ZN(new_n2080_));
  AOI21_X1  g1888(.A(new_n2074_), .B1(new_n2073_), .B2(new_n2079_), .ZN(new_n2081_));
  OAI21_X1  g1889(.A(new_n1976_), .B1(new_n2080_), .B2(new_n2081_), .ZN(new_n2082_));
  INV_X1    g1890(.A(new_n2074_), .ZN(new_n2083_));
  INV_X1    g1891(.A(new_n2079_), .ZN(new_n2084_));
  AOI21_X1  g1892(.A(new_n2075_), .B1(new_n2078_), .B2(new_n1980_), .ZN(new_n2085_));
  OAI21_X1  g1893(.A(new_n2083_), .B1(new_n2084_), .B2(new_n2085_), .ZN(new_n2086_));
  OAI21_X1  g1894(.A(new_n1927_), .B1(new_n1924_), .B2(new_n1810_), .ZN(new_n2087_));
  NAND3_X1  g1895(.A1(new_n2073_), .A2(new_n2074_), .A3(new_n2079_), .ZN(new_n2088_));
  NAND3_X1  g1896(.A1(new_n2086_), .A2(new_n2087_), .A3(new_n2088_), .ZN(new_n2089_));
  NOR2_X1   g1897(.A1(new_n312_), .A2(new_n1405_), .ZN(new_n2090_));
  INV_X1    g1898(.A(new_n2090_), .ZN(new_n2091_));
  AND3_X1   g1899(.A1(new_n2082_), .A2(new_n2089_), .A3(new_n2091_), .ZN(new_n2092_));
  AOI21_X1  g1900(.A(new_n2091_), .B1(new_n2082_), .B2(new_n2089_), .ZN(new_n2093_));
  OAI21_X1  g1901(.A(new_n1975_), .B1(new_n2092_), .B2(new_n2093_), .ZN(new_n2094_));
  NAND2_X1  g1902(.A1(G69gat), .A2(G511gat), .ZN(new_n2095_));
  NOR3_X1   g1903(.A1(new_n2080_), .A2(new_n2081_), .A3(new_n1976_), .ZN(new_n2096_));
  AOI21_X1  g1904(.A(new_n2087_), .B1(new_n2086_), .B2(new_n2088_), .ZN(new_n2097_));
  OAI21_X1  g1905(.A(new_n2090_), .B1(new_n2096_), .B2(new_n2097_), .ZN(new_n2098_));
  NAND3_X1  g1906(.A1(new_n2082_), .A2(new_n2089_), .A3(new_n2091_), .ZN(new_n2099_));
  OAI21_X1  g1907(.A(new_n1935_), .B1(new_n1938_), .B2(new_n1932_), .ZN(new_n2100_));
  NAND3_X1  g1908(.A1(new_n2098_), .A2(new_n2099_), .A3(new_n2100_), .ZN(new_n2101_));
  AND3_X1   g1909(.A1(new_n2094_), .A2(new_n2095_), .A3(new_n2101_), .ZN(new_n2102_));
  AOI21_X1  g1910(.A(new_n2095_), .B1(new_n2094_), .B2(new_n2101_), .ZN(new_n2103_));
  NOR2_X1   g1911(.A1(new_n2102_), .A2(new_n2103_), .ZN(new_n2104_));
  NAND3_X1  g1912(.A1(new_n1941_), .A2(new_n1936_), .A3(new_n1939_), .ZN(new_n2105_));
  NAND2_X1  g1913(.A1(new_n1953_), .A2(new_n2105_), .ZN(new_n2106_));
  NAND2_X1  g1914(.A1(new_n2104_), .A2(new_n2106_), .ZN(new_n2107_));
  NOR2_X1   g1915(.A1(new_n214_), .A2(new_n1622_), .ZN(new_n2108_));
  INV_X1    g1916(.A(new_n2108_), .ZN(new_n2109_));
  OAI211_X1 g1917(.A(new_n1953_), .B(new_n2105_), .C1(new_n2102_), .C2(new_n2103_), .ZN(new_n2110_));
  AND3_X1   g1918(.A1(new_n2107_), .A2(new_n2109_), .A3(new_n2110_), .ZN(new_n2111_));
  AOI21_X1  g1919(.A(new_n2109_), .B1(new_n2107_), .B2(new_n2110_), .ZN(new_n2112_));
  OAI211_X1 g1920(.A(new_n1973_), .B(new_n1974_), .C1(new_n2111_), .C2(new_n2112_), .ZN(new_n2113_));
  NAND2_X1  g1921(.A1(new_n1954_), .A2(new_n1957_), .ZN(new_n2114_));
  NAND2_X1  g1922(.A1(new_n2114_), .A2(new_n1949_), .ZN(new_n2115_));
  NAND2_X1  g1923(.A1(new_n2107_), .A2(new_n2110_), .ZN(new_n2116_));
  NAND2_X1  g1924(.A1(new_n2116_), .A2(new_n2108_), .ZN(new_n2117_));
  NAND3_X1  g1925(.A1(new_n2107_), .A2(new_n2109_), .A3(new_n2110_), .ZN(new_n2118_));
  NAND3_X1  g1926(.A1(new_n2115_), .A2(new_n2117_), .A3(new_n2118_), .ZN(new_n2119_));
  NAND2_X1  g1927(.A1(new_n2113_), .A2(new_n2119_), .ZN(new_n2120_));
  NAND2_X1  g1928(.A1(new_n2117_), .A2(new_n2118_), .ZN(new_n2121_));
  AOI21_X1  g1929(.A(new_n1974_), .B1(new_n2121_), .B2(new_n1973_), .ZN(new_n2122_));
  NOR2_X1   g1930(.A1(new_n2120_), .A2(new_n2122_), .ZN(new_n2123_));
  XNOR2_X1  g1931(.A(new_n1971_), .B(new_n2123_), .ZN(G6170gat));
  OR2_X1    g1932(.A1(new_n2121_), .A2(new_n2115_), .ZN(new_n2125_));
  OAI21_X1  g1933(.A(new_n2125_), .B1(new_n1971_), .B2(new_n2123_), .ZN(new_n2126_));
  NOR2_X1   g1934(.A1(new_n318_), .A2(new_n1622_), .ZN(new_n2127_));
  NOR2_X1   g1935(.A1(new_n2092_), .A2(new_n2096_), .ZN(new_n2128_));
  INV_X1    g1936(.A(new_n2128_), .ZN(new_n2129_));
  AOI21_X1  g1937(.A(new_n2028_), .B1(new_n2033_), .B2(new_n2034_), .ZN(new_n2130_));
  INV_X1    g1938(.A(new_n2130_), .ZN(new_n2131_));
  NOR2_X1   g1939(.A1(new_n1092_), .A2(new_n616_), .ZN(new_n2132_));
  NAND2_X1  g1940(.A1(new_n2024_), .A2(new_n2025_), .ZN(new_n2133_));
  AOI22_X1  g1941(.A1(new_n2133_), .A2(new_n1991_), .B1(new_n2013_), .B2(new_n2017_), .ZN(new_n2134_));
  OR2_X1    g1942(.A1(new_n2011_), .A2(new_n2012_), .ZN(new_n2135_));
  OR2_X1    g1943(.A1(new_n2009_), .A2(new_n2010_), .ZN(new_n2136_));
  NAND2_X1  g1944(.A1(new_n2135_), .A2(new_n2136_), .ZN(new_n2137_));
  NAND3_X1  g1945(.A1(new_n1997_), .A2(new_n2000_), .A3(new_n1998_), .ZN(new_n2138_));
  AND2_X1   g1946(.A1(new_n2138_), .A2(new_n1998_), .ZN(new_n2139_));
  NAND2_X1  g1947(.A1(G256gat), .A2(G341gat), .ZN(new_n2140_));
  XNOR2_X1  g1948(.A(new_n2139_), .B(new_n2140_), .ZN(new_n2141_));
  NAND2_X1  g1949(.A1(new_n348_), .A2(G239gat), .ZN(new_n2142_));
  XOR2_X1   g1950(.A(new_n2141_), .B(new_n2142_), .Z(new_n2143_));
  NOR2_X1   g1951(.A1(new_n1994_), .A2(new_n2001_), .ZN(new_n2144_));
  OAI21_X1  g1952(.A(new_n2002_), .B1(new_n2144_), .B2(new_n2008_), .ZN(new_n2145_));
  XNOR2_X1  g1953(.A(new_n2143_), .B(new_n2145_), .ZN(new_n2146_));
  NAND2_X1  g1954(.A1(G222gat), .A2(G375gat), .ZN(new_n2147_));
  NAND2_X1  g1955(.A1(new_n2146_), .A2(new_n2147_), .ZN(new_n2148_));
  OR2_X1    g1956(.A1(new_n2146_), .A2(new_n2147_), .ZN(new_n2149_));
  NAND3_X1  g1957(.A1(new_n2137_), .A2(new_n2148_), .A3(new_n2149_), .ZN(new_n2150_));
  NAND2_X1  g1958(.A1(new_n2149_), .A2(new_n2148_), .ZN(new_n2151_));
  NAND3_X1  g1959(.A1(new_n2135_), .A2(new_n2136_), .A3(new_n2151_), .ZN(new_n2152_));
  NAND2_X1  g1960(.A1(new_n2150_), .A2(new_n2152_), .ZN(new_n2153_));
  NOR2_X1   g1961(.A1(new_n942_), .A2(new_n867_), .ZN(new_n2154_));
  XNOR2_X1  g1962(.A(new_n2153_), .B(new_n2154_), .ZN(new_n2155_));
  NAND2_X1  g1963(.A1(new_n2134_), .A2(new_n2155_), .ZN(new_n2156_));
  INV_X1    g1964(.A(new_n2156_), .ZN(new_n2157_));
  NOR2_X1   g1965(.A1(new_n2134_), .A2(new_n2155_), .ZN(new_n2158_));
  OAI21_X1  g1966(.A(new_n2132_), .B1(new_n2157_), .B2(new_n2158_), .ZN(new_n2159_));
  INV_X1    g1967(.A(new_n2158_), .ZN(new_n2160_));
  INV_X1    g1968(.A(new_n2132_), .ZN(new_n2161_));
  NAND3_X1  g1969(.A1(new_n2160_), .A2(new_n2161_), .A3(new_n2156_), .ZN(new_n2162_));
  AOI21_X1  g1970(.A(new_n2131_), .B1(new_n2159_), .B2(new_n2162_), .ZN(new_n2163_));
  INV_X1    g1971(.A(new_n2163_), .ZN(new_n2164_));
  NOR2_X1   g1972(.A1(new_n946_), .A2(new_n774_), .ZN(new_n2165_));
  INV_X1    g1973(.A(new_n2165_), .ZN(new_n2166_));
  NAND3_X1  g1974(.A1(new_n2162_), .A2(new_n2131_), .A3(new_n2159_), .ZN(new_n2167_));
  NAND3_X1  g1975(.A1(new_n2164_), .A2(new_n2166_), .A3(new_n2167_), .ZN(new_n2168_));
  INV_X1    g1976(.A(new_n2167_), .ZN(new_n2169_));
  OAI21_X1  g1977(.A(new_n2165_), .B1(new_n2169_), .B2(new_n2163_), .ZN(new_n2170_));
  NAND2_X1  g1978(.A1(new_n2168_), .A2(new_n2170_), .ZN(new_n2171_));
  XNOR2_X1  g1979(.A(new_n2042_), .B(KEYINPUT89), .ZN(new_n2172_));
  NAND3_X1  g1980(.A1(new_n2171_), .A2(new_n2046_), .A3(new_n2172_), .ZN(new_n2173_));
  NAND2_X1  g1981(.A1(new_n2172_), .A2(new_n2046_), .ZN(new_n2174_));
  NAND3_X1  g1982(.A1(new_n2174_), .A2(new_n2168_), .A3(new_n2170_), .ZN(new_n2175_));
  NAND2_X1  g1983(.A1(G154gat), .A2(G443gat), .ZN(new_n2176_));
  NAND3_X1  g1984(.A1(new_n2173_), .A2(new_n2175_), .A3(new_n2176_), .ZN(new_n2177_));
  INV_X1    g1985(.A(new_n2177_), .ZN(new_n2178_));
  AOI21_X1  g1986(.A(new_n2176_), .B1(new_n2173_), .B2(new_n2175_), .ZN(new_n2179_));
  OAI211_X1 g1987(.A(new_n2056_), .B(new_n2057_), .C1(new_n2178_), .C2(new_n2179_), .ZN(new_n2180_));
  INV_X1    g1988(.A(new_n2179_), .ZN(new_n2181_));
  NAND2_X1  g1989(.A1(new_n2057_), .A2(new_n2056_), .ZN(new_n2182_));
  NAND3_X1  g1990(.A1(new_n2181_), .A2(new_n2182_), .A3(new_n2177_), .ZN(new_n2183_));
  NAND2_X1  g1991(.A1(new_n2180_), .A2(new_n2183_), .ZN(new_n2184_));
  NOR2_X1   g1992(.A1(new_n648_), .A2(new_n1055_), .ZN(new_n2185_));
  NAND2_X1  g1993(.A1(new_n2184_), .A2(new_n2185_), .ZN(new_n2186_));
  OAI211_X1 g1994(.A(new_n2180_), .B(new_n2183_), .C1(new_n648_), .C2(new_n1055_), .ZN(new_n2187_));
  NAND2_X1  g1995(.A1(new_n2186_), .A2(new_n2187_), .ZN(new_n2188_));
  NOR2_X1   g1996(.A1(new_n2062_), .A2(new_n2060_), .ZN(new_n2189_));
  OR2_X1    g1997(.A1(new_n2188_), .A2(new_n2189_), .ZN(new_n2190_));
  NAND2_X1  g1998(.A1(new_n2188_), .A2(new_n2189_), .ZN(new_n2191_));
  OR3_X1    g1999(.A1(new_n539_), .A2(new_n1215_), .A3(KEYINPUT90), .ZN(new_n2192_));
  OAI21_X1  g2000(.A(KEYINPUT90), .B1(new_n539_), .B2(new_n1215_), .ZN(new_n2193_));
  AOI22_X1  g2001(.A1(new_n2190_), .A2(new_n2191_), .B1(new_n2192_), .B2(new_n2193_), .ZN(new_n2194_));
  AND2_X1   g2002(.A1(new_n2190_), .A2(new_n2191_), .ZN(new_n2195_));
  AOI21_X1  g2003(.A(new_n2194_), .B1(new_n2195_), .B2(new_n2193_), .ZN(new_n2196_));
  NOR2_X1   g2004(.A1(new_n1978_), .A2(new_n2078_), .ZN(new_n2197_));
  NOR2_X1   g2005(.A1(new_n2081_), .A2(new_n2197_), .ZN(new_n2198_));
  OR2_X1    g2006(.A1(new_n2196_), .A2(new_n2198_), .ZN(new_n2199_));
  NAND2_X1  g2007(.A1(new_n2196_), .A2(new_n2198_), .ZN(new_n2200_));
  NAND2_X1  g2008(.A1(G103gat), .A2(G494gat), .ZN(new_n2201_));
  NAND2_X1  g2009(.A1(new_n2201_), .A2(KEYINPUT91), .ZN(new_n2202_));
  NAND3_X1  g2010(.A1(new_n2199_), .A2(new_n2200_), .A3(new_n2202_), .ZN(new_n2203_));
  INV_X1    g2011(.A(new_n2203_), .ZN(new_n2204_));
  OR2_X1    g2012(.A1(new_n2201_), .A2(KEYINPUT91), .ZN(new_n2205_));
  AOI22_X1  g2013(.A1(new_n2199_), .A2(new_n2200_), .B1(new_n2205_), .B2(new_n2202_), .ZN(new_n2206_));
  OAI21_X1  g2014(.A(new_n2129_), .B1(new_n2204_), .B2(new_n2206_), .ZN(new_n2207_));
  NOR2_X1   g2015(.A1(new_n312_), .A2(new_n1417_), .ZN(new_n2208_));
  INV_X1    g2016(.A(new_n2208_), .ZN(new_n2209_));
  NAND2_X1  g2017(.A1(new_n2199_), .A2(new_n2200_), .ZN(new_n2210_));
  NAND2_X1  g2018(.A1(new_n2205_), .A2(new_n2202_), .ZN(new_n2211_));
  NAND2_X1  g2019(.A1(new_n2210_), .A2(new_n2211_), .ZN(new_n2212_));
  NAND3_X1  g2020(.A1(new_n2212_), .A2(new_n2128_), .A3(new_n2203_), .ZN(new_n2213_));
  NAND3_X1  g2021(.A1(new_n2207_), .A2(new_n2209_), .A3(new_n2213_), .ZN(new_n2214_));
  INV_X1    g2022(.A(new_n2214_), .ZN(new_n2215_));
  INV_X1    g2023(.A(new_n2102_), .ZN(new_n2216_));
  AND2_X1   g2024(.A1(new_n2216_), .A2(new_n2101_), .ZN(new_n2217_));
  AOI21_X1  g2025(.A(new_n2209_), .B1(new_n2207_), .B2(new_n2213_), .ZN(new_n2218_));
  NOR3_X1   g2026(.A1(new_n2215_), .A2(new_n2217_), .A3(new_n2218_), .ZN(new_n2219_));
  NAND2_X1  g2027(.A1(new_n2216_), .A2(new_n2101_), .ZN(new_n2220_));
  INV_X1    g2028(.A(new_n2213_), .ZN(new_n2221_));
  AOI21_X1  g2029(.A(new_n2128_), .B1(new_n2212_), .B2(new_n2203_), .ZN(new_n2222_));
  OAI21_X1  g2030(.A(new_n2208_), .B1(new_n2221_), .B2(new_n2222_), .ZN(new_n2223_));
  AOI21_X1  g2031(.A(new_n2220_), .B1(new_n2223_), .B2(new_n2214_), .ZN(new_n2224_));
  OAI21_X1  g2032(.A(new_n2127_), .B1(new_n2219_), .B2(new_n2224_), .ZN(new_n2225_));
  OAI21_X1  g2033(.A(new_n2217_), .B1(new_n2215_), .B2(new_n2218_), .ZN(new_n2226_));
  NAND3_X1  g2034(.A1(new_n2223_), .A2(new_n2214_), .A3(new_n2220_), .ZN(new_n2227_));
  OAI211_X1 g2035(.A(new_n2226_), .B(new_n2227_), .C1(new_n318_), .C2(new_n1622_), .ZN(new_n2228_));
  NAND2_X1  g2036(.A1(new_n2225_), .A2(new_n2228_), .ZN(new_n2229_));
  NAND2_X1  g2037(.A1(new_n2118_), .A2(new_n2107_), .ZN(new_n2230_));
  XNOR2_X1  g2038(.A(new_n2229_), .B(new_n2230_), .ZN(new_n2231_));
  XNOR2_X1  g2039(.A(new_n2126_), .B(new_n2231_), .ZN(G6180gat));
  AOI21_X1  g2040(.A(new_n2169_), .B1(new_n2164_), .B2(new_n2166_), .ZN(new_n2233_));
  INV_X1    g2041(.A(new_n2233_), .ZN(new_n2234_));
  NAND2_X1  g2042(.A1(G188gat), .A2(G426gat), .ZN(new_n2235_));
  OR2_X1    g2043(.A1(new_n2153_), .A2(new_n2154_), .ZN(new_n2236_));
  NAND2_X1  g2044(.A1(new_n2236_), .A2(new_n2150_), .ZN(new_n2237_));
  OAI211_X1 g2045(.A(new_n2143_), .B(new_n2002_), .C1(new_n2008_), .C2(new_n2144_), .ZN(new_n2238_));
  NAND2_X1  g2046(.A1(new_n2148_), .A2(new_n2238_), .ZN(new_n2239_));
  INV_X1    g2047(.A(KEYINPUT92), .ZN(new_n2240_));
  AOI21_X1  g2048(.A(new_n2240_), .B1(new_n2141_), .B2(new_n2142_), .ZN(new_n2241_));
  INV_X1    g2049(.A(new_n2241_), .ZN(new_n2242_));
  INV_X1    g2050(.A(new_n2139_), .ZN(new_n2243_));
  NAND2_X1  g2051(.A1(new_n2243_), .A2(new_n2140_), .ZN(new_n2244_));
  NAND3_X1  g2052(.A1(new_n2141_), .A2(new_n2240_), .A3(new_n2142_), .ZN(new_n2245_));
  NAND3_X1  g2053(.A1(new_n2242_), .A2(new_n2244_), .A3(new_n2245_), .ZN(new_n2246_));
  OR3_X1    g2054(.A1(new_n2246_), .A2(new_n1823_), .A3(new_n302_), .ZN(new_n2247_));
  NOR2_X1   g2055(.A1(new_n1657_), .A2(new_n356_), .ZN(new_n2248_));
  INV_X1    g2056(.A(new_n2248_), .ZN(new_n2249_));
  OAI21_X1  g2057(.A(new_n2246_), .B1(new_n1823_), .B2(new_n302_), .ZN(new_n2250_));
  NAND3_X1  g2058(.A1(new_n2247_), .A2(new_n2249_), .A3(new_n2250_), .ZN(new_n2251_));
  INV_X1    g2059(.A(new_n2251_), .ZN(new_n2252_));
  AOI21_X1  g2060(.A(new_n2249_), .B1(new_n2247_), .B2(new_n2250_), .ZN(new_n2253_));
  INV_X1    g2061(.A(KEYINPUT93), .ZN(new_n2254_));
  NOR3_X1   g2062(.A1(new_n2252_), .A2(new_n2253_), .A3(new_n2254_), .ZN(new_n2255_));
  NAND2_X1  g2063(.A1(new_n2247_), .A2(new_n2250_), .ZN(new_n2256_));
  NAND2_X1  g2064(.A1(new_n2256_), .A2(new_n2248_), .ZN(new_n2257_));
  AOI21_X1  g2065(.A(KEYINPUT93), .B1(new_n2257_), .B2(new_n2251_), .ZN(new_n2258_));
  OAI21_X1  g2066(.A(new_n2239_), .B1(new_n2255_), .B2(new_n2258_), .ZN(new_n2259_));
  OAI21_X1  g2067(.A(new_n2254_), .B1(new_n2252_), .B2(new_n2253_), .ZN(new_n2260_));
  NAND3_X1  g2068(.A1(new_n2257_), .A2(KEYINPUT93), .A3(new_n2251_), .ZN(new_n2261_));
  NAND4_X1  g2069(.A1(new_n2260_), .A2(new_n2261_), .A3(new_n2238_), .A4(new_n2148_), .ZN(new_n2262_));
  NOR2_X1   g2070(.A1(new_n1437_), .A2(new_n867_), .ZN(new_n2263_));
  INV_X1    g2071(.A(new_n2263_), .ZN(new_n2264_));
  NAND3_X1  g2072(.A1(new_n2259_), .A2(new_n2262_), .A3(new_n2264_), .ZN(new_n2265_));
  NAND2_X1  g2073(.A1(new_n2259_), .A2(new_n2262_), .ZN(new_n2266_));
  NAND2_X1  g2074(.A1(new_n2266_), .A2(new_n2263_), .ZN(new_n2267_));
  NAND3_X1  g2075(.A1(new_n2237_), .A2(new_n2265_), .A3(new_n2267_), .ZN(new_n2268_));
  NAND2_X1  g2076(.A1(new_n2267_), .A2(new_n2265_), .ZN(new_n2269_));
  NAND3_X1  g2077(.A1(new_n2236_), .A2(new_n2269_), .A3(new_n2150_), .ZN(new_n2270_));
  NAND2_X1  g2078(.A1(new_n2268_), .A2(new_n2270_), .ZN(new_n2271_));
  NAND2_X1  g2079(.A1(G205gat), .A2(G409gat), .ZN(new_n2272_));
  XNOR2_X1  g2080(.A(new_n2271_), .B(new_n2272_), .ZN(new_n2273_));
  OAI211_X1 g2081(.A(new_n2160_), .B(KEYINPUT94), .C1(new_n2157_), .C2(new_n2132_), .ZN(new_n2274_));
  OAI21_X1  g2082(.A(new_n2160_), .B1(new_n2157_), .B2(new_n2132_), .ZN(new_n2275_));
  INV_X1    g2083(.A(KEYINPUT94), .ZN(new_n2276_));
  NAND2_X1  g2084(.A1(new_n2275_), .A2(new_n2276_), .ZN(new_n2277_));
  AOI21_X1  g2085(.A(new_n2273_), .B1(new_n2274_), .B2(new_n2277_), .ZN(new_n2278_));
  AND2_X1   g2086(.A1(new_n2273_), .A2(new_n2277_), .ZN(new_n2279_));
  OAI21_X1  g2087(.A(new_n2235_), .B1(new_n2278_), .B2(new_n2279_), .ZN(new_n2280_));
  INV_X1    g2088(.A(new_n2273_), .ZN(new_n2281_));
  NAND2_X1  g2089(.A1(new_n2277_), .A2(new_n2274_), .ZN(new_n2282_));
  NAND2_X1  g2090(.A1(new_n2281_), .A2(new_n2282_), .ZN(new_n2283_));
  NAND2_X1  g2091(.A1(new_n2273_), .A2(new_n2277_), .ZN(new_n2284_));
  NAND4_X1  g2092(.A1(new_n2283_), .A2(G188gat), .A3(G426gat), .A4(new_n2284_), .ZN(new_n2285_));
  AOI21_X1  g2093(.A(new_n2234_), .B1(new_n2280_), .B2(new_n2285_), .ZN(new_n2286_));
  INV_X1    g2094(.A(new_n2286_), .ZN(new_n2287_));
  NOR2_X1   g2095(.A1(new_n946_), .A2(new_n765_), .ZN(new_n2288_));
  INV_X1    g2096(.A(new_n2288_), .ZN(new_n2289_));
  NAND3_X1  g2097(.A1(new_n2280_), .A2(new_n2285_), .A3(new_n2234_), .ZN(new_n2290_));
  NAND3_X1  g2098(.A1(new_n2287_), .A2(new_n2289_), .A3(new_n2290_), .ZN(new_n2291_));
  INV_X1    g2099(.A(new_n2290_), .ZN(new_n2292_));
  OAI21_X1  g2100(.A(new_n2288_), .B1(new_n2292_), .B2(new_n2286_), .ZN(new_n2293_));
  NAND2_X1  g2101(.A1(new_n2291_), .A2(new_n2293_), .ZN(new_n2294_));
  NAND3_X1  g2102(.A1(new_n2294_), .A2(new_n2175_), .A3(new_n2177_), .ZN(new_n2295_));
  NAND2_X1  g2103(.A1(new_n2177_), .A2(new_n2175_), .ZN(new_n2296_));
  NAND3_X1  g2104(.A1(new_n2291_), .A2(new_n2293_), .A3(new_n2296_), .ZN(new_n2297_));
  NAND2_X1  g2105(.A1(new_n2295_), .A2(new_n2297_), .ZN(new_n2298_));
  NAND2_X1  g2106(.A1(G154gat), .A2(G460gat), .ZN(new_n2299_));
  XNOR2_X1  g2107(.A(new_n2299_), .B(KEYINPUT95), .ZN(new_n2300_));
  NAND2_X1  g2108(.A1(new_n2298_), .A2(new_n2300_), .ZN(new_n2301_));
  NAND2_X1  g2109(.A1(new_n2299_), .A2(KEYINPUT95), .ZN(new_n2302_));
  NAND3_X1  g2110(.A1(new_n2295_), .A2(new_n2297_), .A3(new_n2302_), .ZN(new_n2303_));
  NAND2_X1  g2111(.A1(new_n2301_), .A2(new_n2303_), .ZN(new_n2304_));
  NAND2_X1  g2112(.A1(new_n2187_), .A2(new_n2183_), .ZN(new_n2305_));
  NAND2_X1  g2113(.A1(new_n2304_), .A2(new_n2305_), .ZN(new_n2306_));
  NAND4_X1  g2114(.A1(new_n2301_), .A2(new_n2183_), .A3(new_n2187_), .A4(new_n2303_), .ZN(new_n2307_));
  NAND2_X1  g2115(.A1(new_n2306_), .A2(new_n2307_), .ZN(new_n2308_));
  NAND3_X1  g2116(.A1(new_n2308_), .A2(G137gat), .A3(G477gat), .ZN(new_n2309_));
  NAND2_X1  g2117(.A1(G137gat), .A2(G477gat), .ZN(new_n2310_));
  XNOR2_X1  g2118(.A(new_n2310_), .B(KEYINPUT96), .ZN(new_n2311_));
  NAND3_X1  g2119(.A1(new_n2306_), .A2(new_n2307_), .A3(new_n2311_), .ZN(new_n2312_));
  NAND2_X1  g2120(.A1(new_n2309_), .A2(new_n2312_), .ZN(new_n2313_));
  INV_X1    g2121(.A(new_n2191_), .ZN(new_n2314_));
  AND3_X1   g2122(.A1(new_n2190_), .A2(G120gat), .A3(G477gat), .ZN(new_n2315_));
  OAI21_X1  g2123(.A(new_n2313_), .B1(new_n2314_), .B2(new_n2315_), .ZN(new_n2316_));
  NAND2_X1  g2124(.A1(G120gat), .A2(G494gat), .ZN(new_n2317_));
  NOR2_X1   g2125(.A1(new_n2315_), .A2(new_n2314_), .ZN(new_n2318_));
  NAND3_X1  g2126(.A1(new_n2318_), .A2(new_n2309_), .A3(new_n2312_), .ZN(new_n2319_));
  AND3_X1   g2127(.A1(new_n2316_), .A2(new_n2317_), .A3(new_n2319_), .ZN(new_n2320_));
  AOI21_X1  g2128(.A(new_n2317_), .B1(new_n2316_), .B2(new_n2319_), .ZN(new_n2321_));
  NOR2_X1   g2129(.A1(new_n2320_), .A2(new_n2321_), .ZN(new_n2322_));
  NAND2_X1  g2130(.A1(new_n2200_), .A2(new_n2201_), .ZN(new_n2323_));
  NAND2_X1  g2131(.A1(new_n2323_), .A2(new_n2199_), .ZN(new_n2324_));
  OR2_X1    g2132(.A1(new_n2322_), .A2(new_n2324_), .ZN(new_n2325_));
  NAND2_X1  g2133(.A1(new_n2322_), .A2(new_n2324_), .ZN(new_n2326_));
  NAND2_X1  g2134(.A1(new_n2325_), .A2(new_n2326_), .ZN(new_n2327_));
  NOR2_X1   g2135(.A1(new_n455_), .A2(new_n1417_), .ZN(new_n2328_));
  NAND2_X1  g2136(.A1(new_n2327_), .A2(new_n2328_), .ZN(new_n2329_));
  INV_X1    g2137(.A(new_n2328_), .ZN(new_n2330_));
  NAND3_X1  g2138(.A1(new_n2325_), .A2(new_n2330_), .A3(new_n2326_), .ZN(new_n2331_));
  NAND2_X1  g2139(.A1(new_n2329_), .A2(new_n2331_), .ZN(new_n2332_));
  NOR2_X1   g2140(.A1(new_n2215_), .A2(new_n2222_), .ZN(new_n2333_));
  XNOR2_X1  g2141(.A(new_n2332_), .B(new_n2333_), .ZN(new_n2334_));
  NAND2_X1  g2142(.A1(G86gat), .A2(G528gat), .ZN(new_n2335_));
  XNOR2_X1  g2143(.A(new_n2334_), .B(new_n2335_), .ZN(new_n2336_));
  NAND2_X1  g2144(.A1(new_n2228_), .A2(new_n2227_), .ZN(new_n2337_));
  NAND2_X1  g2145(.A1(new_n2336_), .A2(new_n2337_), .ZN(new_n2338_));
  INV_X1    g2146(.A(new_n2338_), .ZN(new_n2339_));
  NOR2_X1   g2147(.A1(new_n2336_), .A2(new_n2337_), .ZN(new_n2340_));
  NOR2_X1   g2148(.A1(new_n2339_), .A2(new_n2340_), .ZN(new_n2341_));
  AOI21_X1  g2149(.A(new_n2229_), .B1(new_n2107_), .B2(new_n2118_), .ZN(new_n2342_));
  AOI21_X1  g2150(.A(new_n2342_), .B1(new_n2126_), .B2(new_n2231_), .ZN(new_n2343_));
  XOR2_X1   g2151(.A(new_n2341_), .B(new_n2343_), .Z(G6190gat));
  OAI21_X1  g2152(.A(new_n2338_), .B1(new_n2343_), .B2(new_n2340_), .ZN(new_n2345_));
  XNOR2_X1  g2153(.A(new_n2345_), .B(KEYINPUT106), .ZN(new_n2346_));
  NOR2_X1   g2154(.A1(new_n455_), .A2(new_n1622_), .ZN(new_n2347_));
  INV_X1    g2155(.A(new_n2319_), .ZN(new_n2348_));
  AOI21_X1  g2156(.A(new_n2348_), .B1(new_n2317_), .B2(new_n2316_), .ZN(new_n2349_));
  INV_X1    g2157(.A(new_n2349_), .ZN(new_n2350_));
  NOR2_X1   g2158(.A1(new_n957_), .A2(new_n1215_), .ZN(new_n2351_));
  INV_X1    g2159(.A(new_n2351_), .ZN(new_n2352_));
  NAND3_X1  g2160(.A1(new_n2297_), .A2(G154gat), .A3(G460gat), .ZN(new_n2353_));
  NAND2_X1  g2161(.A1(new_n2353_), .A2(new_n2295_), .ZN(new_n2354_));
  INV_X1    g2162(.A(KEYINPUT101), .ZN(new_n2355_));
  NOR2_X1   g2163(.A1(new_n946_), .A2(new_n1055_), .ZN(new_n2356_));
  INV_X1    g2164(.A(new_n2356_), .ZN(new_n2357_));
  NOR2_X1   g2165(.A1(new_n1092_), .A2(new_n765_), .ZN(new_n2358_));
  AOI21_X1  g2166(.A(KEYINPUT98), .B1(new_n2265_), .B2(new_n2259_), .ZN(new_n2359_));
  INV_X1    g2167(.A(new_n2359_), .ZN(new_n2360_));
  NOR2_X1   g2168(.A1(new_n1823_), .A2(new_n356_), .ZN(new_n2361_));
  XNOR2_X1  g2169(.A(new_n2361_), .B(KEYINPUT97), .ZN(new_n2362_));
  NAND3_X1  g2170(.A1(new_n2251_), .A2(new_n2250_), .A3(new_n2362_), .ZN(new_n2363_));
  INV_X1    g2171(.A(new_n2363_), .ZN(new_n2364_));
  NAND2_X1  g2172(.A1(new_n2251_), .A2(new_n2250_), .ZN(new_n2365_));
  AOI21_X1  g2173(.A(new_n2364_), .B1(new_n2361_), .B2(new_n2365_), .ZN(new_n2366_));
  NOR2_X1   g2174(.A1(new_n1657_), .A2(new_n867_), .ZN(new_n2367_));
  AND2_X1   g2175(.A1(new_n2366_), .A2(new_n2367_), .ZN(new_n2368_));
  NOR2_X1   g2176(.A1(new_n2366_), .A2(new_n2367_), .ZN(new_n2369_));
  NOR2_X1   g2177(.A1(new_n2368_), .A2(new_n2369_), .ZN(new_n2370_));
  INV_X1    g2178(.A(new_n2370_), .ZN(new_n2371_));
  NOR3_X1   g2179(.A1(new_n2255_), .A2(new_n2258_), .A3(new_n2239_), .ZN(new_n2372_));
  OAI211_X1 g2180(.A(KEYINPUT98), .B(new_n2259_), .C1(new_n2372_), .C2(new_n2263_), .ZN(new_n2373_));
  NAND3_X1  g2181(.A1(new_n2360_), .A2(new_n2371_), .A3(new_n2373_), .ZN(new_n2374_));
  INV_X1    g2182(.A(new_n2373_), .ZN(new_n2375_));
  OAI21_X1  g2183(.A(new_n2370_), .B1(new_n2375_), .B2(new_n2359_), .ZN(new_n2376_));
  NOR2_X1   g2184(.A1(new_n1437_), .A2(new_n616_), .ZN(new_n2377_));
  INV_X1    g2185(.A(new_n2377_), .ZN(new_n2378_));
  AND3_X1   g2186(.A1(new_n2374_), .A2(new_n2376_), .A3(new_n2378_), .ZN(new_n2379_));
  AOI21_X1  g2187(.A(new_n2378_), .B1(new_n2374_), .B2(new_n2376_), .ZN(new_n2380_));
  NOR2_X1   g2188(.A1(new_n2379_), .A2(new_n2380_), .ZN(new_n2381_));
  NAND3_X1  g2189(.A1(new_n2268_), .A2(new_n2272_), .A3(new_n2270_), .ZN(new_n2382_));
  NAND2_X1  g2190(.A1(new_n2382_), .A2(new_n2268_), .ZN(new_n2383_));
  NAND2_X1  g2191(.A1(new_n2381_), .A2(new_n2383_), .ZN(new_n2384_));
  OAI211_X1 g2192(.A(new_n2382_), .B(new_n2268_), .C1(new_n2379_), .C2(new_n2380_), .ZN(new_n2385_));
  NAND2_X1  g2193(.A1(new_n2384_), .A2(new_n2385_), .ZN(new_n2386_));
  NAND3_X1  g2194(.A1(new_n2386_), .A2(G205gat), .A3(G426gat), .ZN(new_n2387_));
  OAI211_X1 g2195(.A(new_n2384_), .B(new_n2385_), .C1(new_n942_), .C2(new_n774_), .ZN(new_n2388_));
  NAND2_X1  g2196(.A1(new_n2387_), .A2(new_n2388_), .ZN(new_n2389_));
  NAND2_X1  g2197(.A1(new_n2273_), .A2(new_n2275_), .ZN(new_n2390_));
  AND3_X1   g2198(.A1(new_n2280_), .A2(new_n2389_), .A3(new_n2390_), .ZN(new_n2391_));
  AOI21_X1  g2199(.A(new_n2389_), .B1(new_n2280_), .B2(new_n2390_), .ZN(new_n2392_));
  OAI21_X1  g2200(.A(new_n2358_), .B1(new_n2391_), .B2(new_n2392_), .ZN(new_n2393_));
  NAND2_X1  g2201(.A1(new_n2280_), .A2(new_n2390_), .ZN(new_n2394_));
  AND2_X1   g2202(.A1(new_n2387_), .A2(new_n2388_), .ZN(new_n2395_));
  NAND2_X1  g2203(.A1(new_n2394_), .A2(new_n2395_), .ZN(new_n2396_));
  INV_X1    g2204(.A(new_n2358_), .ZN(new_n2397_));
  NAND3_X1  g2205(.A1(new_n2280_), .A2(new_n2389_), .A3(new_n2390_), .ZN(new_n2398_));
  NAND3_X1  g2206(.A1(new_n2396_), .A2(new_n2397_), .A3(new_n2398_), .ZN(new_n2399_));
  NAND2_X1  g2207(.A1(new_n2393_), .A2(new_n2399_), .ZN(new_n2400_));
  OAI21_X1  g2208(.A(new_n2290_), .B1(new_n2286_), .B2(new_n2288_), .ZN(new_n2401_));
  INV_X1    g2209(.A(KEYINPUT99), .ZN(new_n2402_));
  NAND2_X1  g2210(.A1(new_n2401_), .A2(new_n2402_), .ZN(new_n2403_));
  OAI211_X1 g2211(.A(KEYINPUT99), .B(new_n2290_), .C1(new_n2286_), .C2(new_n2288_), .ZN(new_n2404_));
  AOI21_X1  g2212(.A(new_n2400_), .B1(new_n2403_), .B2(new_n2404_), .ZN(new_n2405_));
  AND2_X1   g2213(.A1(new_n2400_), .A2(new_n2404_), .ZN(new_n2406_));
  OAI21_X1  g2214(.A(new_n2357_), .B1(new_n2405_), .B2(new_n2406_), .ZN(new_n2407_));
  INV_X1    g2215(.A(new_n2400_), .ZN(new_n2408_));
  NAND2_X1  g2216(.A1(new_n2403_), .A2(new_n2404_), .ZN(new_n2409_));
  NAND2_X1  g2217(.A1(new_n2408_), .A2(new_n2409_), .ZN(new_n2410_));
  NAND2_X1  g2218(.A1(new_n2400_), .A2(new_n2404_), .ZN(new_n2411_));
  NAND3_X1  g2219(.A1(new_n2410_), .A2(new_n2356_), .A3(new_n2411_), .ZN(new_n2412_));
  AND3_X1   g2220(.A1(new_n2407_), .A2(KEYINPUT100), .A3(new_n2412_), .ZN(new_n2413_));
  AOI21_X1  g2221(.A(KEYINPUT100), .B1(new_n2407_), .B2(new_n2412_), .ZN(new_n2414_));
  OAI21_X1  g2222(.A(new_n2355_), .B1(new_n2413_), .B2(new_n2414_), .ZN(new_n2415_));
  INV_X1    g2223(.A(KEYINPUT100), .ZN(new_n2416_));
  NOR3_X1   g2224(.A1(new_n2405_), .A2(new_n2406_), .A3(new_n2357_), .ZN(new_n2417_));
  AOI21_X1  g2225(.A(new_n2356_), .B1(new_n2410_), .B2(new_n2411_), .ZN(new_n2418_));
  OAI21_X1  g2226(.A(new_n2416_), .B1(new_n2417_), .B2(new_n2418_), .ZN(new_n2419_));
  NAND3_X1  g2227(.A1(new_n2407_), .A2(new_n2412_), .A3(KEYINPUT100), .ZN(new_n2420_));
  NAND3_X1  g2228(.A1(new_n2419_), .A2(KEYINPUT101), .A3(new_n2420_), .ZN(new_n2421_));
  AOI21_X1  g2229(.A(new_n2354_), .B1(new_n2415_), .B2(new_n2421_), .ZN(new_n2422_));
  INV_X1    g2230(.A(new_n2354_), .ZN(new_n2423_));
  NAND2_X1  g2231(.A1(new_n2419_), .A2(new_n2420_), .ZN(new_n2424_));
  AOI21_X1  g2232(.A(new_n2423_), .B1(new_n2424_), .B2(new_n2355_), .ZN(new_n2425_));
  OAI21_X1  g2233(.A(new_n2352_), .B1(new_n2422_), .B2(new_n2425_), .ZN(new_n2426_));
  NOR3_X1   g2234(.A1(new_n2413_), .A2(new_n2414_), .A3(new_n2355_), .ZN(new_n2427_));
  AOI21_X1  g2235(.A(KEYINPUT101), .B1(new_n2419_), .B2(new_n2420_), .ZN(new_n2428_));
  OAI21_X1  g2236(.A(new_n2423_), .B1(new_n2427_), .B2(new_n2428_), .ZN(new_n2429_));
  NAND2_X1  g2237(.A1(new_n2415_), .A2(new_n2354_), .ZN(new_n2430_));
  NAND3_X1  g2238(.A1(new_n2429_), .A2(new_n2351_), .A3(new_n2430_), .ZN(new_n2431_));
  NAND2_X1  g2239(.A1(new_n2312_), .A2(new_n2306_), .ZN(new_n2432_));
  AND3_X1   g2240(.A1(new_n2426_), .A2(new_n2431_), .A3(new_n2432_), .ZN(new_n2433_));
  AOI21_X1  g2241(.A(new_n2432_), .B1(new_n2426_), .B2(new_n2431_), .ZN(new_n2434_));
  NOR2_X1   g2242(.A1(new_n648_), .A2(new_n1405_), .ZN(new_n2435_));
  NOR3_X1   g2243(.A1(new_n2433_), .A2(new_n2434_), .A3(new_n2435_), .ZN(new_n2436_));
  INV_X1    g2244(.A(new_n2435_), .ZN(new_n2437_));
  INV_X1    g2245(.A(new_n2432_), .ZN(new_n2438_));
  AOI21_X1  g2246(.A(new_n2351_), .B1(new_n2429_), .B2(new_n2430_), .ZN(new_n2439_));
  NOR3_X1   g2247(.A1(new_n2422_), .A2(new_n2352_), .A3(new_n2425_), .ZN(new_n2440_));
  OAI21_X1  g2248(.A(new_n2438_), .B1(new_n2439_), .B2(new_n2440_), .ZN(new_n2441_));
  NAND3_X1  g2249(.A1(new_n2426_), .A2(new_n2431_), .A3(new_n2432_), .ZN(new_n2442_));
  AOI21_X1  g2250(.A(new_n2437_), .B1(new_n2441_), .B2(new_n2442_), .ZN(new_n2443_));
  OAI21_X1  g2251(.A(new_n2350_), .B1(new_n2436_), .B2(new_n2443_), .ZN(new_n2444_));
  INV_X1    g2252(.A(KEYINPUT103), .ZN(new_n2445_));
  NAND2_X1  g2253(.A1(new_n2444_), .A2(new_n2445_), .ZN(new_n2446_));
  OAI21_X1  g2254(.A(new_n2435_), .B1(new_n2433_), .B2(new_n2434_), .ZN(new_n2447_));
  NAND3_X1  g2255(.A1(new_n2441_), .A2(new_n2437_), .A3(new_n2442_), .ZN(new_n2448_));
  NAND2_X1  g2256(.A1(new_n2447_), .A2(new_n2448_), .ZN(new_n2449_));
  NAND3_X1  g2257(.A1(new_n2449_), .A2(KEYINPUT103), .A3(new_n2350_), .ZN(new_n2450_));
  NAND2_X1  g2258(.A1(new_n2446_), .A2(new_n2450_), .ZN(new_n2451_));
  NOR2_X1   g2259(.A1(new_n539_), .A2(new_n1417_), .ZN(new_n2452_));
  NAND3_X1  g2260(.A1(new_n2447_), .A2(new_n2349_), .A3(new_n2448_), .ZN(new_n2453_));
  NAND2_X1  g2261(.A1(new_n2453_), .A2(KEYINPUT102), .ZN(new_n2454_));
  INV_X1    g2262(.A(KEYINPUT102), .ZN(new_n2455_));
  NAND4_X1  g2263(.A1(new_n2447_), .A2(new_n2448_), .A3(new_n2455_), .A4(new_n2349_), .ZN(new_n2456_));
  NAND2_X1  g2264(.A1(new_n2454_), .A2(new_n2456_), .ZN(new_n2457_));
  AND3_X1   g2265(.A1(new_n2451_), .A2(new_n2452_), .A3(new_n2457_), .ZN(new_n2458_));
  AOI21_X1  g2266(.A(new_n2452_), .B1(new_n2451_), .B2(new_n2457_), .ZN(new_n2459_));
  NAND2_X1  g2267(.A1(new_n2331_), .A2(new_n2326_), .ZN(new_n2460_));
  INV_X1    g2268(.A(new_n2460_), .ZN(new_n2461_));
  NOR3_X1   g2269(.A1(new_n2458_), .A2(new_n2459_), .A3(new_n2461_), .ZN(new_n2462_));
  AOI21_X1  g2270(.A(KEYINPUT103), .B1(new_n2449_), .B2(new_n2350_), .ZN(new_n2463_));
  AOI211_X1 g2271(.A(new_n2445_), .B(new_n2349_), .C1(new_n2447_), .C2(new_n2448_), .ZN(new_n2464_));
  OAI21_X1  g2272(.A(new_n2457_), .B1(new_n2463_), .B2(new_n2464_), .ZN(new_n2465_));
  INV_X1    g2273(.A(new_n2452_), .ZN(new_n2466_));
  NAND2_X1  g2274(.A1(new_n2465_), .A2(new_n2466_), .ZN(new_n2467_));
  NAND3_X1  g2275(.A1(new_n2451_), .A2(new_n2452_), .A3(new_n2457_), .ZN(new_n2468_));
  AOI21_X1  g2276(.A(new_n2460_), .B1(new_n2467_), .B2(new_n2468_), .ZN(new_n2469_));
  OAI21_X1  g2277(.A(new_n2347_), .B1(new_n2462_), .B2(new_n2469_), .ZN(new_n2470_));
  OAI21_X1  g2278(.A(new_n2461_), .B1(new_n2458_), .B2(new_n2459_), .ZN(new_n2471_));
  NAND3_X1  g2279(.A1(new_n2467_), .A2(new_n2460_), .A3(new_n2468_), .ZN(new_n2472_));
  INV_X1    g2280(.A(new_n2347_), .ZN(new_n2473_));
  NAND3_X1  g2281(.A1(new_n2471_), .A2(new_n2472_), .A3(new_n2473_), .ZN(new_n2474_));
  NOR2_X1   g2282(.A1(new_n2332_), .A2(new_n2333_), .ZN(new_n2475_));
  NAND2_X1  g2283(.A1(new_n2332_), .A2(new_n2333_), .ZN(new_n2476_));
  AOI21_X1  g2284(.A(new_n2475_), .B1(new_n2335_), .B2(new_n2476_), .ZN(new_n2477_));
  NAND3_X1  g2285(.A1(new_n2470_), .A2(new_n2474_), .A3(new_n2477_), .ZN(new_n2478_));
  INV_X1    g2286(.A(KEYINPUT105), .ZN(new_n2479_));
  NAND2_X1  g2287(.A1(new_n2478_), .A2(new_n2479_), .ZN(new_n2480_));
  NAND4_X1  g2288(.A1(new_n2470_), .A2(KEYINPUT105), .A3(new_n2474_), .A4(new_n2477_), .ZN(new_n2481_));
  NAND2_X1  g2289(.A1(new_n2480_), .A2(new_n2481_), .ZN(new_n2482_));
  INV_X1    g2290(.A(new_n2477_), .ZN(new_n2483_));
  OAI21_X1  g2291(.A(KEYINPUT104), .B1(new_n2462_), .B2(new_n2469_), .ZN(new_n2484_));
  NAND2_X1  g2292(.A1(new_n2470_), .A2(new_n2474_), .ZN(new_n2485_));
  OAI211_X1 g2293(.A(new_n2483_), .B(new_n2484_), .C1(new_n2485_), .C2(KEYINPUT104), .ZN(new_n2486_));
  NAND2_X1  g2294(.A1(new_n2482_), .A2(new_n2486_), .ZN(new_n2487_));
  XNOR2_X1  g2295(.A(new_n2346_), .B(new_n2487_), .ZN(G6200gat));
  NOR2_X1   g2296(.A1(new_n2485_), .A2(new_n2477_), .ZN(new_n2489_));
  AOI21_X1  g2297(.A(new_n2489_), .B1(new_n2345_), .B2(new_n2487_), .ZN(new_n2490_));
  NAND2_X1  g2298(.A1(new_n2474_), .A2(new_n2472_), .ZN(new_n2491_));
  INV_X1    g2299(.A(new_n2491_), .ZN(new_n2492_));
  INV_X1    g2300(.A(KEYINPUT109), .ZN(new_n2493_));
  NAND2_X1  g2301(.A1(new_n2365_), .A2(new_n2362_), .ZN(new_n2494_));
  OAI21_X1  g2302(.A(new_n2494_), .B1(new_n2366_), .B2(new_n2367_), .ZN(new_n2495_));
  NAND2_X1  g2303(.A1(G256gat), .A2(G392gat), .ZN(new_n2496_));
  XNOR2_X1  g2304(.A(new_n2495_), .B(new_n2496_), .ZN(new_n2497_));
  NOR2_X1   g2305(.A1(new_n1657_), .A2(new_n616_), .ZN(new_n2498_));
  OR2_X1    g2306(.A1(new_n2497_), .A2(new_n2498_), .ZN(new_n2499_));
  NAND2_X1  g2307(.A1(new_n2497_), .A2(new_n2498_), .ZN(new_n2500_));
  INV_X1    g2308(.A(KEYINPUT107), .ZN(new_n2501_));
  OAI21_X1  g2309(.A(new_n2376_), .B1(new_n2379_), .B2(new_n2501_), .ZN(new_n2502_));
  NAND3_X1  g2310(.A1(new_n2374_), .A2(new_n2376_), .A3(new_n2378_), .ZN(new_n2503_));
  NOR2_X1   g2311(.A1(new_n2503_), .A2(KEYINPUT107), .ZN(new_n2504_));
  OAI211_X1 g2312(.A(new_n2499_), .B(new_n2500_), .C1(new_n2502_), .C2(new_n2504_), .ZN(new_n2505_));
  NAND2_X1  g2313(.A1(new_n2499_), .A2(new_n2500_), .ZN(new_n2506_));
  NAND3_X1  g2314(.A1(new_n2506_), .A2(new_n2376_), .A3(new_n2503_), .ZN(new_n2507_));
  NAND2_X1  g2315(.A1(new_n2505_), .A2(new_n2507_), .ZN(new_n2508_));
  NAND3_X1  g2316(.A1(new_n2508_), .A2(G222gat), .A3(G426gat), .ZN(new_n2509_));
  OAI211_X1 g2317(.A(new_n2505_), .B(new_n2507_), .C1(new_n1437_), .C2(new_n774_), .ZN(new_n2510_));
  AND2_X1   g2318(.A1(new_n2509_), .A2(new_n2510_), .ZN(new_n2511_));
  NAND2_X1  g2319(.A1(new_n2388_), .A2(new_n2384_), .ZN(new_n2512_));
  OR2_X1    g2320(.A1(new_n2511_), .A2(new_n2512_), .ZN(new_n2513_));
  NAND2_X1  g2321(.A1(new_n2511_), .A2(new_n2512_), .ZN(new_n2514_));
  AND2_X1   g2322(.A1(new_n2513_), .A2(new_n2514_), .ZN(new_n2515_));
  NOR2_X1   g2323(.A1(new_n942_), .A2(new_n765_), .ZN(new_n2516_));
  XNOR2_X1  g2324(.A(new_n2516_), .B(KEYINPUT108), .ZN(new_n2517_));
  AND2_X1   g2325(.A1(new_n2515_), .A2(new_n2517_), .ZN(new_n2518_));
  AND2_X1   g2326(.A1(new_n2516_), .A2(KEYINPUT108), .ZN(new_n2519_));
  NOR2_X1   g2327(.A1(new_n2515_), .A2(new_n2519_), .ZN(new_n2520_));
  OAI21_X1  g2328(.A(new_n2493_), .B1(new_n2518_), .B2(new_n2520_), .ZN(new_n2521_));
  NAND2_X1  g2329(.A1(new_n2515_), .A2(new_n2517_), .ZN(new_n2522_));
  OAI211_X1 g2330(.A(new_n2522_), .B(KEYINPUT109), .C1(new_n2515_), .C2(new_n2519_), .ZN(new_n2523_));
  AND2_X1   g2331(.A1(new_n2521_), .A2(new_n2523_), .ZN(new_n2524_));
  NAND2_X1  g2332(.A1(new_n2399_), .A2(new_n2396_), .ZN(new_n2525_));
  NAND2_X1  g2333(.A1(new_n2524_), .A2(new_n2525_), .ZN(new_n2526_));
  NOR2_X1   g2334(.A1(new_n1092_), .A2(new_n1055_), .ZN(new_n2527_));
  INV_X1    g2335(.A(new_n2527_), .ZN(new_n2528_));
  INV_X1    g2336(.A(new_n2525_), .ZN(new_n2529_));
  OAI211_X1 g2337(.A(new_n2522_), .B(new_n2529_), .C1(new_n2515_), .C2(new_n2519_), .ZN(new_n2530_));
  NAND3_X1  g2338(.A1(new_n2526_), .A2(new_n2528_), .A3(new_n2530_), .ZN(new_n2531_));
  NAND2_X1  g2339(.A1(new_n2521_), .A2(new_n2523_), .ZN(new_n2532_));
  OAI21_X1  g2340(.A(new_n2530_), .B1(new_n2532_), .B2(new_n2529_), .ZN(new_n2533_));
  NAND2_X1  g2341(.A1(new_n2533_), .A2(new_n2527_), .ZN(new_n2534_));
  AND3_X1   g2342(.A1(new_n2531_), .A2(KEYINPUT110), .A3(new_n2534_), .ZN(new_n2535_));
  AOI21_X1  g2343(.A(KEYINPUT110), .B1(new_n2531_), .B2(new_n2534_), .ZN(new_n2536_));
  NOR2_X1   g2344(.A1(new_n2535_), .A2(new_n2536_), .ZN(new_n2537_));
  AOI21_X1  g2345(.A(new_n2400_), .B1(new_n2290_), .B2(new_n2291_), .ZN(new_n2538_));
  OR2_X1    g2346(.A1(new_n2418_), .A2(new_n2538_), .ZN(new_n2539_));
  NOR2_X1   g2347(.A1(new_n946_), .A2(new_n1215_), .ZN(new_n2540_));
  XOR2_X1   g2348(.A(new_n2539_), .B(new_n2540_), .Z(new_n2541_));
  NAND2_X1  g2349(.A1(new_n2537_), .A2(new_n2541_), .ZN(new_n2542_));
  NAND2_X1  g2350(.A1(new_n2531_), .A2(new_n2534_), .ZN(new_n2543_));
  OAI21_X1  g2351(.A(new_n2542_), .B1(new_n2543_), .B2(new_n2541_), .ZN(new_n2544_));
  NOR2_X1   g2352(.A1(new_n2424_), .A2(new_n2354_), .ZN(new_n2545_));
  NOR2_X1   g2353(.A1(new_n2439_), .A2(new_n2545_), .ZN(new_n2546_));
  AND2_X1   g2354(.A1(new_n2544_), .A2(new_n2546_), .ZN(new_n2547_));
  NOR2_X1   g2355(.A1(new_n2544_), .A2(new_n2546_), .ZN(new_n2548_));
  OAI211_X1 g2356(.A(G154gat), .B(G494gat), .C1(new_n2547_), .C2(new_n2548_), .ZN(new_n2549_));
  INV_X1    g2357(.A(new_n2548_), .ZN(new_n2550_));
  NAND2_X1  g2358(.A1(G154gat), .A2(G494gat), .ZN(new_n2551_));
  NAND2_X1  g2359(.A1(new_n2544_), .A2(new_n2546_), .ZN(new_n2552_));
  NAND3_X1  g2360(.A1(new_n2550_), .A2(new_n2551_), .A3(new_n2552_), .ZN(new_n2553_));
  AND2_X1   g2361(.A1(new_n2549_), .A2(new_n2553_), .ZN(new_n2554_));
  NAND2_X1  g2362(.A1(new_n2448_), .A2(new_n2442_), .ZN(new_n2555_));
  XNOR2_X1  g2363(.A(new_n2555_), .B(KEYINPUT111), .ZN(new_n2556_));
  NAND2_X1  g2364(.A1(new_n2554_), .A2(new_n2556_), .ZN(new_n2557_));
  NAND2_X1  g2365(.A1(new_n2549_), .A2(new_n2553_), .ZN(new_n2558_));
  OAI21_X1  g2366(.A(new_n2558_), .B1(KEYINPUT111), .B2(new_n2555_), .ZN(new_n2559_));
  NAND2_X1  g2367(.A1(new_n2557_), .A2(new_n2559_), .ZN(new_n2560_));
  NAND2_X1  g2368(.A1(G137gat), .A2(G511gat), .ZN(new_n2561_));
  NAND2_X1  g2369(.A1(new_n2560_), .A2(new_n2561_), .ZN(new_n2562_));
  NAND4_X1  g2370(.A1(new_n2557_), .A2(new_n2559_), .A3(G137gat), .A4(G511gat), .ZN(new_n2563_));
  NAND2_X1  g2371(.A1(new_n2562_), .A2(new_n2563_), .ZN(new_n2564_));
  NAND3_X1  g2372(.A1(new_n2350_), .A2(new_n2447_), .A3(new_n2448_), .ZN(new_n2565_));
  NAND3_X1  g2373(.A1(new_n2564_), .A2(new_n2467_), .A3(new_n2565_), .ZN(new_n2566_));
  NOR2_X1   g2374(.A1(new_n539_), .A2(new_n1622_), .ZN(new_n2567_));
  INV_X1    g2375(.A(new_n2567_), .ZN(new_n2568_));
  NAND2_X1  g2376(.A1(new_n2467_), .A2(new_n2565_), .ZN(new_n2569_));
  NAND3_X1  g2377(.A1(new_n2562_), .A2(new_n2569_), .A3(new_n2563_), .ZN(new_n2570_));
  NAND3_X1  g2378(.A1(new_n2566_), .A2(new_n2568_), .A3(new_n2570_), .ZN(new_n2571_));
  INV_X1    g2379(.A(new_n2571_), .ZN(new_n2572_));
  AOI21_X1  g2380(.A(new_n2568_), .B1(new_n2566_), .B2(new_n2570_), .ZN(new_n2573_));
  OAI21_X1  g2381(.A(new_n2492_), .B1(new_n2572_), .B2(new_n2573_), .ZN(new_n2574_));
  INV_X1    g2382(.A(new_n2573_), .ZN(new_n2575_));
  NAND3_X1  g2383(.A1(new_n2575_), .A2(new_n2491_), .A3(new_n2571_), .ZN(new_n2576_));
  NAND2_X1  g2384(.A1(new_n2574_), .A2(new_n2576_), .ZN(new_n2577_));
  XNOR2_X1  g2385(.A(new_n2490_), .B(new_n2577_), .ZN(G6210gat));
  OAI21_X1  g2386(.A(new_n2576_), .B1(new_n2490_), .B2(new_n2577_), .ZN(new_n2579_));
  INV_X1    g2387(.A(new_n2539_), .ZN(new_n2580_));
  OAI21_X1  g2388(.A(new_n2580_), .B1(new_n2537_), .B2(new_n2540_), .ZN(new_n2581_));
  NAND2_X1  g2389(.A1(new_n2543_), .A2(new_n2540_), .ZN(new_n2582_));
  NAND2_X1  g2390(.A1(new_n2581_), .A2(new_n2582_), .ZN(new_n2583_));
  AOI22_X1  g2391(.A1(new_n2524_), .A2(new_n2525_), .B1(new_n2528_), .B2(new_n2530_), .ZN(new_n2584_));
  INV_X1    g2392(.A(new_n2584_), .ZN(new_n2585_));
  NAND2_X1  g2393(.A1(new_n2514_), .A2(new_n2516_), .ZN(new_n2586_));
  NAND2_X1  g2394(.A1(new_n2586_), .A2(new_n2513_), .ZN(new_n2587_));
  XNOR2_X1  g2395(.A(new_n2587_), .B(KEYINPUT114), .ZN(new_n2588_));
  NOR2_X1   g2396(.A1(new_n1657_), .A2(new_n774_), .ZN(new_n2589_));
  INV_X1    g2397(.A(new_n2589_), .ZN(new_n2590_));
  OAI21_X1  g2398(.A(new_n2495_), .B1(new_n1823_), .B2(new_n867_), .ZN(new_n2591_));
  NAND2_X1  g2399(.A1(new_n2499_), .A2(new_n2591_), .ZN(new_n2592_));
  OAI21_X1  g2400(.A(new_n2592_), .B1(new_n1823_), .B2(new_n616_), .ZN(new_n2593_));
  NAND4_X1  g2401(.A1(new_n2499_), .A2(G256gat), .A3(G409gat), .A4(new_n2591_), .ZN(new_n2594_));
  AOI21_X1  g2402(.A(new_n2590_), .B1(new_n2593_), .B2(new_n2594_), .ZN(new_n2595_));
  INV_X1    g2403(.A(new_n2595_), .ZN(new_n2596_));
  NAND3_X1  g2404(.A1(new_n2593_), .A2(new_n2590_), .A3(new_n2594_), .ZN(new_n2597_));
  NAND2_X1  g2405(.A1(new_n2596_), .A2(new_n2597_), .ZN(new_n2598_));
  XNOR2_X1  g2406(.A(new_n2598_), .B(KEYINPUT113), .ZN(new_n2599_));
  XNOR2_X1  g2407(.A(new_n2505_), .B(KEYINPUT112), .ZN(new_n2600_));
  NAND2_X1  g2408(.A1(new_n2600_), .A2(new_n2510_), .ZN(new_n2601_));
  NOR2_X1   g2409(.A1(new_n2599_), .A2(new_n2601_), .ZN(new_n2602_));
  NAND3_X1  g2410(.A1(new_n2596_), .A2(KEYINPUT113), .A3(new_n2597_), .ZN(new_n2603_));
  AND2_X1   g2411(.A1(new_n2601_), .A2(new_n2603_), .ZN(new_n2604_));
  NOR2_X1   g2412(.A1(new_n2602_), .A2(new_n2604_), .ZN(new_n2605_));
  NAND3_X1  g2413(.A1(new_n2605_), .A2(G222gat), .A3(G443gat), .ZN(new_n2606_));
  OAI22_X1  g2414(.A1(new_n2602_), .A2(new_n2604_), .B1(new_n1437_), .B2(new_n765_), .ZN(new_n2607_));
  NAND3_X1  g2415(.A1(new_n2588_), .A2(new_n2606_), .A3(new_n2607_), .ZN(new_n2608_));
  NOR2_X1   g2416(.A1(new_n942_), .A2(new_n1055_), .ZN(new_n2609_));
  INV_X1    g2417(.A(new_n2609_), .ZN(new_n2610_));
  NAND2_X1  g2418(.A1(new_n2606_), .A2(new_n2607_), .ZN(new_n2611_));
  NAND2_X1  g2419(.A1(new_n2611_), .A2(new_n2587_), .ZN(new_n2612_));
  NAND3_X1  g2420(.A1(new_n2608_), .A2(new_n2610_), .A3(new_n2612_), .ZN(new_n2613_));
  INV_X1    g2421(.A(new_n2613_), .ZN(new_n2614_));
  AOI21_X1  g2422(.A(new_n2610_), .B1(new_n2608_), .B2(new_n2612_), .ZN(new_n2615_));
  OAI21_X1  g2423(.A(new_n2585_), .B1(new_n2614_), .B2(new_n2615_), .ZN(new_n2616_));
  INV_X1    g2424(.A(KEYINPUT115), .ZN(new_n2617_));
  NOR2_X1   g2425(.A1(new_n2614_), .A2(new_n2615_), .ZN(new_n2618_));
  NAND2_X1  g2426(.A1(new_n2618_), .A2(new_n2584_), .ZN(new_n2619_));
  NAND3_X1  g2427(.A1(new_n2616_), .A2(new_n2617_), .A3(new_n2619_), .ZN(new_n2620_));
  NAND3_X1  g2428(.A1(new_n2618_), .A2(KEYINPUT115), .A3(new_n2584_), .ZN(new_n2621_));
  NOR2_X1   g2429(.A1(new_n1092_), .A2(new_n1215_), .ZN(new_n2622_));
  INV_X1    g2430(.A(new_n2622_), .ZN(new_n2623_));
  NAND3_X1  g2431(.A1(new_n2620_), .A2(new_n2621_), .A3(new_n2623_), .ZN(new_n2624_));
  NAND2_X1  g2432(.A1(new_n2616_), .A2(new_n2619_), .ZN(new_n2625_));
  OAI21_X1  g2433(.A(new_n2624_), .B1(new_n2623_), .B2(new_n2625_), .ZN(new_n2626_));
  NAND2_X1  g2434(.A1(new_n2583_), .A2(new_n2626_), .ZN(new_n2627_));
  NOR2_X1   g2435(.A1(new_n946_), .A2(new_n1405_), .ZN(new_n2628_));
  INV_X1    g2436(.A(new_n2628_), .ZN(new_n2629_));
  NAND2_X1  g2437(.A1(new_n2620_), .A2(new_n2621_), .ZN(new_n2630_));
  NAND2_X1  g2438(.A1(new_n2630_), .A2(new_n2622_), .ZN(new_n2631_));
  NAND2_X1  g2439(.A1(new_n2625_), .A2(new_n2623_), .ZN(new_n2632_));
  NAND4_X1  g2440(.A1(new_n2631_), .A2(new_n2581_), .A3(new_n2582_), .A4(new_n2632_), .ZN(new_n2633_));
  NAND3_X1  g2441(.A1(new_n2627_), .A2(new_n2629_), .A3(new_n2633_), .ZN(new_n2634_));
  INV_X1    g2442(.A(new_n2634_), .ZN(new_n2635_));
  AOI21_X1  g2443(.A(new_n2629_), .B1(new_n2627_), .B2(new_n2633_), .ZN(new_n2636_));
  NOR2_X1   g2444(.A1(new_n2635_), .A2(new_n2636_), .ZN(new_n2637_));
  NAND2_X1  g2445(.A1(new_n2553_), .A2(new_n2550_), .ZN(new_n2638_));
  NAND2_X1  g2446(.A1(new_n2637_), .A2(new_n2638_), .ZN(new_n2639_));
  OAI211_X1 g2447(.A(new_n2553_), .B(new_n2550_), .C1(new_n2635_), .C2(new_n2636_), .ZN(new_n2640_));
  NAND2_X1  g2448(.A1(new_n2639_), .A2(new_n2640_), .ZN(new_n2641_));
  NOR2_X1   g2449(.A1(new_n957_), .A2(new_n1417_), .ZN(new_n2642_));
  INV_X1    g2450(.A(new_n2642_), .ZN(new_n2643_));
  XNOR2_X1  g2451(.A(new_n2641_), .B(new_n2643_), .ZN(new_n2644_));
  NAND2_X1  g2452(.A1(new_n2554_), .A2(new_n2555_), .ZN(new_n2645_));
  NAND2_X1  g2453(.A1(new_n2562_), .A2(new_n2645_), .ZN(new_n2646_));
  NAND2_X1  g2454(.A1(new_n2644_), .A2(new_n2646_), .ZN(new_n2647_));
  INV_X1    g2455(.A(new_n2647_), .ZN(new_n2648_));
  NOR2_X1   g2456(.A1(new_n2644_), .A2(new_n2646_), .ZN(new_n2649_));
  OAI211_X1 g2457(.A(G137gat), .B(G528gat), .C1(new_n2648_), .C2(new_n2649_), .ZN(new_n2650_));
  INV_X1    g2458(.A(new_n2649_), .ZN(new_n2651_));
  NAND2_X1  g2459(.A1(G137gat), .A2(G528gat), .ZN(new_n2652_));
  NAND3_X1  g2460(.A1(new_n2651_), .A2(new_n2652_), .A3(new_n2647_), .ZN(new_n2653_));
  NAND2_X1  g2461(.A1(new_n2650_), .A2(new_n2653_), .ZN(new_n2654_));
  NAND2_X1  g2462(.A1(new_n2571_), .A2(new_n2570_), .ZN(new_n2655_));
  XNOR2_X1  g2463(.A(new_n2654_), .B(new_n2655_), .ZN(new_n2656_));
  XNOR2_X1  g2464(.A(new_n2579_), .B(new_n2656_), .ZN(G6220gat));
  AOI21_X1  g2465(.A(new_n2654_), .B1(new_n2570_), .B2(new_n2571_), .ZN(new_n2658_));
  AOI21_X1  g2466(.A(new_n2658_), .B1(new_n2579_), .B2(new_n2656_), .ZN(new_n2659_));
  NAND2_X1  g2467(.A1(new_n2585_), .A2(new_n2618_), .ZN(new_n2660_));
  NAND2_X1  g2468(.A1(new_n2624_), .A2(new_n2660_), .ZN(new_n2661_));
  NAND2_X1  g2469(.A1(new_n2613_), .A2(new_n2608_), .ZN(new_n2662_));
  NAND2_X1  g2470(.A1(new_n2597_), .A2(new_n2593_), .ZN(new_n2663_));
  XNOR2_X1  g2471(.A(new_n2663_), .B(KEYINPUT117), .ZN(new_n2664_));
  AOI21_X1  g2472(.A(new_n2664_), .B1(G256gat), .B2(G426gat), .ZN(new_n2665_));
  INV_X1    g2473(.A(new_n2665_), .ZN(new_n2666_));
  NAND3_X1  g2474(.A1(new_n2664_), .A2(G256gat), .A3(G426gat), .ZN(new_n2667_));
  NAND2_X1  g2475(.A1(new_n2666_), .A2(new_n2667_), .ZN(new_n2668_));
  NOR2_X1   g2476(.A1(new_n1657_), .A2(new_n765_), .ZN(new_n2669_));
  INV_X1    g2477(.A(new_n2669_), .ZN(new_n2670_));
  XNOR2_X1  g2478(.A(new_n2668_), .B(new_n2670_), .ZN(new_n2671_));
  INV_X1    g2479(.A(new_n2601_), .ZN(new_n2672_));
  OAI21_X1  g2480(.A(new_n2607_), .B1(new_n2672_), .B2(new_n2598_), .ZN(new_n2673_));
  XNOR2_X1  g2481(.A(new_n2671_), .B(new_n2673_), .ZN(new_n2674_));
  NOR2_X1   g2482(.A1(new_n1437_), .A2(new_n1055_), .ZN(new_n2675_));
  OR2_X1    g2483(.A1(new_n2674_), .A2(new_n2675_), .ZN(new_n2676_));
  NAND2_X1  g2484(.A1(new_n2674_), .A2(new_n2675_), .ZN(new_n2677_));
  AOI21_X1  g2485(.A(new_n2662_), .B1(new_n2676_), .B2(new_n2677_), .ZN(new_n2678_));
  INV_X1    g2486(.A(new_n2678_), .ZN(new_n2679_));
  NAND3_X1  g2487(.A1(new_n2676_), .A2(new_n2677_), .A3(new_n2662_), .ZN(new_n2680_));
  OAI211_X1 g2488(.A(new_n2679_), .B(new_n2680_), .C1(new_n942_), .C2(new_n1215_), .ZN(new_n2681_));
  NAND2_X1  g2489(.A1(new_n2679_), .A2(new_n2680_), .ZN(new_n2682_));
  NOR2_X1   g2490(.A1(new_n942_), .A2(new_n1215_), .ZN(new_n2683_));
  NAND2_X1  g2491(.A1(new_n2682_), .A2(new_n2683_), .ZN(new_n2684_));
  NAND3_X1  g2492(.A1(new_n2661_), .A2(new_n2681_), .A3(new_n2684_), .ZN(new_n2685_));
  NAND2_X1  g2493(.A1(new_n2684_), .A2(new_n2681_), .ZN(new_n2686_));
  NAND3_X1  g2494(.A1(new_n2686_), .A2(new_n2632_), .A3(new_n2660_), .ZN(new_n2687_));
  NAND2_X1  g2495(.A1(new_n2685_), .A2(new_n2687_), .ZN(new_n2688_));
  NOR2_X1   g2496(.A1(new_n1092_), .A2(new_n1405_), .ZN(new_n2689_));
  NAND2_X1  g2497(.A1(new_n2688_), .A2(new_n2689_), .ZN(new_n2690_));
  INV_X1    g2498(.A(new_n2689_), .ZN(new_n2691_));
  NAND3_X1  g2499(.A1(new_n2685_), .A2(new_n2691_), .A3(new_n2687_), .ZN(new_n2692_));
  NAND2_X1  g2500(.A1(new_n2690_), .A2(new_n2692_), .ZN(new_n2693_));
  OR2_X1    g2501(.A1(new_n2693_), .A2(KEYINPUT118), .ZN(new_n2694_));
  NAND2_X1  g2502(.A1(new_n2693_), .A2(KEYINPUT118), .ZN(new_n2695_));
  OR2_X1    g2503(.A1(new_n2634_), .A2(KEYINPUT116), .ZN(new_n2696_));
  NOR2_X1   g2504(.A1(new_n2583_), .A2(new_n2626_), .ZN(new_n2697_));
  AOI21_X1  g2505(.A(new_n2697_), .B1(new_n2634_), .B2(KEYINPUT116), .ZN(new_n2698_));
  NAND2_X1  g2506(.A1(new_n2696_), .A2(new_n2698_), .ZN(new_n2699_));
  NAND3_X1  g2507(.A1(new_n2694_), .A2(new_n2695_), .A3(new_n2699_), .ZN(new_n2700_));
  NAND4_X1  g2508(.A1(new_n2696_), .A2(new_n2698_), .A3(new_n2693_), .A4(KEYINPUT118), .ZN(new_n2701_));
  NAND2_X1  g2509(.A1(new_n2700_), .A2(new_n2701_), .ZN(new_n2702_));
  NOR2_X1   g2510(.A1(new_n946_), .A2(new_n1417_), .ZN(new_n2703_));
  NAND2_X1  g2511(.A1(new_n2702_), .A2(new_n2703_), .ZN(new_n2704_));
  INV_X1    g2512(.A(new_n2703_), .ZN(new_n2705_));
  NAND3_X1  g2513(.A1(new_n2700_), .A2(new_n2705_), .A3(new_n2701_), .ZN(new_n2706_));
  NAND2_X1  g2514(.A1(new_n2704_), .A2(new_n2706_), .ZN(new_n2707_));
  NAND2_X1  g2515(.A1(new_n2707_), .A2(KEYINPUT119), .ZN(new_n2708_));
  INV_X1    g2516(.A(KEYINPUT119), .ZN(new_n2709_));
  NAND3_X1  g2517(.A1(new_n2704_), .A2(new_n2709_), .A3(new_n2706_), .ZN(new_n2710_));
  NAND3_X1  g2518(.A1(new_n2639_), .A2(new_n2643_), .A3(new_n2640_), .ZN(new_n2711_));
  NAND2_X1  g2519(.A1(new_n2711_), .A2(new_n2639_), .ZN(new_n2712_));
  NAND3_X1  g2520(.A1(new_n2708_), .A2(new_n2710_), .A3(new_n2712_), .ZN(new_n2713_));
  AOI21_X1  g2521(.A(new_n2712_), .B1(new_n2704_), .B2(new_n2706_), .ZN(new_n2714_));
  INV_X1    g2522(.A(new_n2714_), .ZN(new_n2715_));
  NAND2_X1  g2523(.A1(new_n2713_), .A2(new_n2715_), .ZN(new_n2716_));
  NOR2_X1   g2524(.A1(new_n957_), .A2(new_n1622_), .ZN(new_n2717_));
  NAND2_X1  g2525(.A1(new_n2716_), .A2(new_n2717_), .ZN(new_n2718_));
  OAI211_X1 g2526(.A(new_n2713_), .B(new_n2715_), .C1(new_n957_), .C2(new_n1622_), .ZN(new_n2719_));
  NAND2_X1  g2527(.A1(new_n2718_), .A2(new_n2719_), .ZN(new_n2720_));
  AOI21_X1  g2528(.A(new_n2648_), .B1(new_n2651_), .B2(new_n2652_), .ZN(new_n2721_));
  NAND2_X1  g2529(.A1(new_n2720_), .A2(new_n2721_), .ZN(new_n2722_));
  INV_X1    g2530(.A(new_n2721_), .ZN(new_n2723_));
  NAND3_X1  g2531(.A1(new_n2718_), .A2(new_n2723_), .A3(new_n2719_), .ZN(new_n2724_));
  NAND2_X1  g2532(.A1(new_n2722_), .A2(new_n2724_), .ZN(new_n2725_));
  XNOR2_X1  g2533(.A(new_n2659_), .B(new_n2725_), .ZN(G6230gat));
  OAI21_X1  g2534(.A(new_n2724_), .B1(new_n2659_), .B2(new_n2725_), .ZN(new_n2727_));
  NAND3_X1  g2535(.A1(new_n2699_), .A2(new_n2692_), .A3(new_n2690_), .ZN(new_n2728_));
  NAND2_X1  g2536(.A1(new_n2706_), .A2(new_n2728_), .ZN(new_n2729_));
  AND2_X1   g2537(.A1(new_n2692_), .A2(new_n2685_), .ZN(new_n2730_));
  NAND2_X1  g2538(.A1(new_n2671_), .A2(new_n2673_), .ZN(new_n2731_));
  OAI21_X1  g2539(.A(new_n2731_), .B1(new_n2674_), .B2(new_n2675_), .ZN(new_n2732_));
  AOI21_X1  g2540(.A(new_n2665_), .B1(new_n2670_), .B2(new_n2667_), .ZN(new_n2733_));
  NOR2_X1   g2541(.A1(new_n1823_), .A2(new_n765_), .ZN(new_n2734_));
  OR2_X1    g2542(.A1(new_n2733_), .A2(new_n2734_), .ZN(new_n2735_));
  NAND2_X1  g2543(.A1(G239gat), .A2(G460gat), .ZN(new_n2736_));
  NAND2_X1  g2544(.A1(new_n2733_), .A2(new_n2734_), .ZN(new_n2737_));
  NAND3_X1  g2545(.A1(new_n2735_), .A2(new_n2736_), .A3(new_n2737_), .ZN(new_n2738_));
  INV_X1    g2546(.A(new_n2738_), .ZN(new_n2739_));
  AOI21_X1  g2547(.A(new_n2736_), .B1(new_n2735_), .B2(new_n2737_), .ZN(new_n2740_));
  NOR2_X1   g2548(.A1(new_n2739_), .A2(new_n2740_), .ZN(new_n2741_));
  OR2_X1    g2549(.A1(new_n2732_), .A2(new_n2741_), .ZN(new_n2742_));
  NAND2_X1  g2550(.A1(new_n2732_), .A2(new_n2741_), .ZN(new_n2743_));
  AOI211_X1 g2551(.A(new_n1437_), .B(new_n1215_), .C1(new_n2742_), .C2(new_n2743_), .ZN(new_n2744_));
  NAND2_X1  g2552(.A1(new_n2742_), .A2(new_n2743_), .ZN(new_n2745_));
  NOR2_X1   g2553(.A1(new_n1437_), .A2(new_n1215_), .ZN(new_n2746_));
  NOR2_X1   g2554(.A1(new_n2745_), .A2(new_n2746_), .ZN(new_n2747_));
  NOR2_X1   g2555(.A1(new_n2744_), .A2(new_n2747_), .ZN(new_n2748_));
  NAND2_X1  g2556(.A1(new_n2681_), .A2(new_n2680_), .ZN(new_n2749_));
  NAND2_X1  g2557(.A1(new_n2748_), .A2(new_n2749_), .ZN(new_n2750_));
  NOR2_X1   g2558(.A1(new_n942_), .A2(new_n1405_), .ZN(new_n2751_));
  INV_X1    g2559(.A(new_n2751_), .ZN(new_n2752_));
  OAI211_X1 g2560(.A(new_n2680_), .B(new_n2681_), .C1(new_n2744_), .C2(new_n2747_), .ZN(new_n2753_));
  AND3_X1   g2561(.A1(new_n2750_), .A2(new_n2752_), .A3(new_n2753_), .ZN(new_n2754_));
  AOI21_X1  g2562(.A(new_n2752_), .B1(new_n2750_), .B2(new_n2753_), .ZN(new_n2755_));
  OR2_X1    g2563(.A1(new_n2754_), .A2(new_n2755_), .ZN(new_n2756_));
  AND2_X1   g2564(.A1(new_n2730_), .A2(new_n2756_), .ZN(new_n2757_));
  NOR2_X1   g2565(.A1(new_n2730_), .A2(new_n2756_), .ZN(new_n2758_));
  NOR2_X1   g2566(.A1(new_n2757_), .A2(new_n2758_), .ZN(new_n2759_));
  OAI21_X1  g2567(.A(new_n2759_), .B1(new_n1092_), .B2(new_n1417_), .ZN(new_n2760_));
  OAI211_X1 g2568(.A(G188gat), .B(G511gat), .C1(new_n2757_), .C2(new_n2758_), .ZN(new_n2761_));
  NAND3_X1  g2569(.A1(new_n2729_), .A2(new_n2760_), .A3(new_n2761_), .ZN(new_n2762_));
  NAND2_X1  g2570(.A1(new_n2760_), .A2(new_n2761_), .ZN(new_n2763_));
  NAND3_X1  g2571(.A1(new_n2763_), .A2(new_n2706_), .A3(new_n2728_), .ZN(new_n2764_));
  NAND2_X1  g2572(.A1(new_n2762_), .A2(new_n2764_), .ZN(new_n2765_));
  NAND3_X1  g2573(.A1(new_n2765_), .A2(G171gat), .A3(G528gat), .ZN(new_n2766_));
  OAI211_X1 g2574(.A(new_n2762_), .B(new_n2764_), .C1(new_n946_), .C2(new_n1622_), .ZN(new_n2767_));
  NAND2_X1  g2575(.A1(new_n2766_), .A2(new_n2767_), .ZN(new_n2768_));
  NAND3_X1  g2576(.A1(new_n2719_), .A2(new_n2768_), .A3(new_n2713_), .ZN(new_n2769_));
  OAI21_X1  g2577(.A(new_n2713_), .B1(new_n2714_), .B2(new_n2717_), .ZN(new_n2770_));
  NAND3_X1  g2578(.A1(new_n2770_), .A2(new_n2766_), .A3(new_n2767_), .ZN(new_n2771_));
  AND3_X1   g2579(.A1(new_n2769_), .A2(new_n2771_), .A3(KEYINPUT120), .ZN(new_n2772_));
  AOI21_X1  g2580(.A(KEYINPUT120), .B1(new_n2769_), .B2(new_n2771_), .ZN(new_n2773_));
  NOR3_X1   g2581(.A1(new_n2772_), .A2(new_n2773_), .A3(KEYINPUT121), .ZN(new_n2774_));
  NOR2_X1   g2582(.A1(new_n2727_), .A2(new_n2774_), .ZN(new_n2775_));
  NOR2_X1   g2583(.A1(new_n2772_), .A2(new_n2773_), .ZN(new_n2776_));
  XOR2_X1   g2584(.A(new_n2776_), .B(KEYINPUT121), .Z(new_n2777_));
  AOI21_X1  g2585(.A(new_n2775_), .B1(new_n2777_), .B2(new_n2727_), .ZN(G6240gat));
  OAI211_X1 g2586(.A(new_n2724_), .B(new_n2771_), .C1(new_n2659_), .C2(new_n2725_), .ZN(new_n2779_));
  NAND2_X1  g2587(.A1(new_n2779_), .A2(new_n2769_), .ZN(new_n2780_));
  INV_X1    g2588(.A(new_n2754_), .ZN(new_n2781_));
  NAND2_X1  g2589(.A1(new_n2781_), .A2(new_n2750_), .ZN(new_n2782_));
  OAI21_X1  g2590(.A(new_n2743_), .B1(new_n2745_), .B2(new_n2746_), .ZN(new_n2783_));
  NAND2_X1  g2591(.A1(new_n2738_), .A2(new_n2735_), .ZN(new_n2784_));
  OAI21_X1  g2592(.A(new_n2784_), .B1(new_n1823_), .B2(new_n1055_), .ZN(new_n2785_));
  NAND4_X1  g2593(.A1(new_n2738_), .A2(G256gat), .A3(G460gat), .A4(new_n2735_), .ZN(new_n2786_));
  NAND2_X1  g2594(.A1(new_n2785_), .A2(new_n2786_), .ZN(new_n2787_));
  NOR2_X1   g2595(.A1(new_n1657_), .A2(new_n1215_), .ZN(new_n2788_));
  XOR2_X1   g2596(.A(new_n2787_), .B(new_n2788_), .Z(new_n2789_));
  OR2_X1    g2597(.A1(new_n2783_), .A2(new_n2789_), .ZN(new_n2790_));
  NAND2_X1  g2598(.A1(new_n2783_), .A2(new_n2789_), .ZN(new_n2791_));
  NAND2_X1  g2599(.A1(new_n2790_), .A2(new_n2791_), .ZN(new_n2792_));
  NAND2_X1  g2600(.A1(G222gat), .A2(G494gat), .ZN(new_n2793_));
  XNOR2_X1  g2601(.A(new_n2792_), .B(new_n2793_), .ZN(new_n2794_));
  OR2_X1    g2602(.A1(new_n2782_), .A2(new_n2794_), .ZN(new_n2795_));
  NAND2_X1  g2603(.A1(new_n2782_), .A2(new_n2794_), .ZN(new_n2796_));
  NAND2_X1  g2604(.A1(new_n2795_), .A2(new_n2796_), .ZN(new_n2797_));
  NAND2_X1  g2605(.A1(G205gat), .A2(G511gat), .ZN(new_n2798_));
  XOR2_X1   g2606(.A(new_n2797_), .B(new_n2798_), .Z(new_n2799_));
  INV_X1    g2607(.A(new_n2758_), .ZN(new_n2800_));
  AND2_X1   g2608(.A1(new_n2760_), .A2(new_n2800_), .ZN(new_n2801_));
  OR2_X1    g2609(.A1(new_n2799_), .A2(new_n2801_), .ZN(new_n2802_));
  NAND2_X1  g2610(.A1(new_n2799_), .A2(new_n2801_), .ZN(new_n2803_));
  NAND2_X1  g2611(.A1(new_n2802_), .A2(new_n2803_), .ZN(new_n2804_));
  NAND2_X1  g2612(.A1(G188gat), .A2(G528gat), .ZN(new_n2805_));
  XNOR2_X1  g2613(.A(new_n2804_), .B(new_n2805_), .ZN(new_n2806_));
  NAND2_X1  g2614(.A1(new_n2767_), .A2(new_n2762_), .ZN(new_n2807_));
  XNOR2_X1  g2615(.A(new_n2806_), .B(new_n2807_), .ZN(new_n2808_));
  NAND2_X1  g2616(.A1(new_n2780_), .A2(new_n2808_), .ZN(new_n2809_));
  INV_X1    g2617(.A(new_n2808_), .ZN(new_n2810_));
  NAND3_X1  g2618(.A1(new_n2779_), .A2(new_n2769_), .A3(new_n2810_), .ZN(new_n2811_));
  NAND2_X1  g2619(.A1(new_n2809_), .A2(new_n2811_), .ZN(G6250gat));
  NAND2_X1  g2620(.A1(new_n2806_), .A2(new_n2807_), .ZN(new_n2813_));
  NAND3_X1  g2621(.A1(new_n2802_), .A2(new_n2805_), .A3(new_n2803_), .ZN(new_n2814_));
  NAND2_X1  g2622(.A1(new_n2814_), .A2(new_n2802_), .ZN(new_n2815_));
  XNOR2_X1  g2623(.A(new_n2815_), .B(KEYINPUT123), .ZN(new_n2816_));
  NAND3_X1  g2624(.A1(new_n2790_), .A2(new_n2793_), .A3(new_n2791_), .ZN(new_n2817_));
  NAND2_X1  g2625(.A1(new_n2817_), .A2(new_n2791_), .ZN(new_n2818_));
  OAI21_X1  g2626(.A(new_n2785_), .B1(new_n2787_), .B2(new_n2788_), .ZN(new_n2819_));
  OR3_X1    g2627(.A1(new_n2819_), .A2(new_n1823_), .A3(new_n1215_), .ZN(new_n2820_));
  OAI21_X1  g2628(.A(new_n2819_), .B1(new_n1823_), .B2(new_n1215_), .ZN(new_n2821_));
  NAND2_X1  g2629(.A1(new_n2820_), .A2(new_n2821_), .ZN(new_n2822_));
  NOR2_X1   g2630(.A1(new_n1657_), .A2(new_n1405_), .ZN(new_n2823_));
  XOR2_X1   g2631(.A(new_n2822_), .B(new_n2823_), .Z(new_n2824_));
  XNOR2_X1  g2632(.A(new_n2818_), .B(new_n2824_), .ZN(new_n2825_));
  XNOR2_X1  g2633(.A(new_n2825_), .B(KEYINPUT122), .ZN(new_n2826_));
  OR3_X1    g2634(.A1(new_n2826_), .A2(new_n1437_), .A3(new_n1417_), .ZN(new_n2827_));
  OAI21_X1  g2635(.A(new_n2826_), .B1(new_n1437_), .B2(new_n1417_), .ZN(new_n2828_));
  NAND2_X1  g2636(.A1(new_n2827_), .A2(new_n2828_), .ZN(new_n2829_));
  NAND3_X1  g2637(.A1(new_n2795_), .A2(new_n2796_), .A3(new_n2798_), .ZN(new_n2830_));
  NAND2_X1  g2638(.A1(new_n2830_), .A2(new_n2796_), .ZN(new_n2831_));
  XNOR2_X1  g2639(.A(new_n2829_), .B(new_n2831_), .ZN(new_n2832_));
  NAND2_X1  g2640(.A1(G205gat), .A2(G528gat), .ZN(new_n2833_));
  XNOR2_X1  g2641(.A(new_n2832_), .B(new_n2833_), .ZN(new_n2834_));
  OR2_X1    g2642(.A1(new_n2816_), .A2(new_n2834_), .ZN(new_n2835_));
  NAND2_X1  g2643(.A1(new_n2816_), .A2(new_n2834_), .ZN(new_n2836_));
  NAND2_X1  g2644(.A1(new_n2835_), .A2(new_n2836_), .ZN(new_n2837_));
  NAND3_X1  g2645(.A1(new_n2811_), .A2(new_n2813_), .A3(new_n2837_), .ZN(new_n2838_));
  AOI21_X1  g2646(.A(new_n2808_), .B1(new_n2776_), .B2(new_n2771_), .ZN(new_n2839_));
  NAND2_X1  g2647(.A1(new_n2779_), .A2(new_n2839_), .ZN(new_n2840_));
  NAND2_X1  g2648(.A1(new_n2840_), .A2(KEYINPUT124), .ZN(new_n2841_));
  INV_X1    g2649(.A(KEYINPUT124), .ZN(new_n2842_));
  NAND3_X1  g2650(.A1(new_n2779_), .A2(new_n2842_), .A3(new_n2839_), .ZN(new_n2843_));
  NAND3_X1  g2651(.A1(new_n2841_), .A2(new_n2813_), .A3(new_n2843_), .ZN(new_n2844_));
  INV_X1    g2652(.A(new_n2844_), .ZN(new_n2845_));
  OAI21_X1  g2653(.A(new_n2838_), .B1(new_n2845_), .B2(new_n2837_), .ZN(G6260gat));
  NAND3_X1  g2654(.A1(new_n2811_), .A2(new_n2813_), .A3(new_n2835_), .ZN(new_n2847_));
  NAND2_X1  g2655(.A1(new_n2847_), .A2(new_n2836_), .ZN(new_n2848_));
  NAND2_X1  g2656(.A1(new_n2818_), .A2(new_n2824_), .ZN(new_n2849_));
  NAND2_X1  g2657(.A1(new_n2828_), .A2(new_n2849_), .ZN(new_n2850_));
  OAI21_X1  g2658(.A(new_n2821_), .B1(new_n2822_), .B2(new_n2823_), .ZN(new_n2851_));
  OR3_X1    g2659(.A1(new_n2851_), .A2(new_n1823_), .A3(new_n1405_), .ZN(new_n2852_));
  OAI21_X1  g2660(.A(new_n2851_), .B1(new_n1823_), .B2(new_n1405_), .ZN(new_n2853_));
  NAND2_X1  g2661(.A1(new_n2852_), .A2(new_n2853_), .ZN(new_n2854_));
  XOR2_X1   g2662(.A(new_n2854_), .B(KEYINPUT125), .Z(new_n2855_));
  NAND2_X1  g2663(.A1(G239gat), .A2(G511gat), .ZN(new_n2856_));
  NAND2_X1  g2664(.A1(new_n2855_), .A2(new_n2856_), .ZN(new_n2857_));
  INV_X1    g2665(.A(new_n2857_), .ZN(new_n2858_));
  NOR2_X1   g2666(.A1(new_n2855_), .A2(new_n2856_), .ZN(new_n2859_));
  NOR2_X1   g2667(.A1(new_n2858_), .A2(new_n2859_), .ZN(new_n2860_));
  XOR2_X1   g2668(.A(new_n2850_), .B(new_n2860_), .Z(new_n2861_));
  OR3_X1    g2669(.A1(new_n2861_), .A2(new_n1437_), .A3(new_n1622_), .ZN(new_n2862_));
  OAI21_X1  g2670(.A(new_n2861_), .B1(new_n1437_), .B2(new_n1622_), .ZN(new_n2863_));
  AND2_X1   g2671(.A1(new_n2862_), .A2(new_n2863_), .ZN(new_n2864_));
  NAND2_X1  g2672(.A1(new_n2832_), .A2(new_n2833_), .ZN(new_n2865_));
  NAND3_X1  g2673(.A1(new_n2827_), .A2(new_n2831_), .A3(new_n2828_), .ZN(new_n2866_));
  NAND2_X1  g2674(.A1(new_n2865_), .A2(new_n2866_), .ZN(new_n2867_));
  NOR2_X1   g2675(.A1(new_n2864_), .A2(new_n2867_), .ZN(new_n2868_));
  INV_X1    g2676(.A(new_n2868_), .ZN(new_n2869_));
  NAND2_X1  g2677(.A1(new_n2864_), .A2(new_n2867_), .ZN(new_n2870_));
  AND2_X1   g2678(.A1(new_n2869_), .A2(new_n2870_), .ZN(new_n2871_));
  XOR2_X1   g2679(.A(new_n2848_), .B(new_n2871_), .Z(G6270gat));
  INV_X1    g2680(.A(KEYINPUT126), .ZN(new_n2873_));
  OAI21_X1  g2681(.A(new_n2853_), .B1(new_n2857_), .B2(new_n2873_), .ZN(new_n2874_));
  AOI21_X1  g2682(.A(new_n2874_), .B1(new_n2873_), .B2(new_n2857_), .ZN(new_n2875_));
  INV_X1    g2683(.A(new_n2875_), .ZN(new_n2876_));
  NOR2_X1   g2684(.A1(new_n1823_), .A2(new_n1417_), .ZN(new_n2877_));
  INV_X1    g2685(.A(new_n2877_), .ZN(new_n2878_));
  NOR2_X1   g2686(.A1(new_n2876_), .A2(new_n2878_), .ZN(new_n2879_));
  INV_X1    g2687(.A(new_n2879_), .ZN(new_n2880_));
  NAND2_X1  g2688(.A1(new_n2876_), .A2(new_n2878_), .ZN(new_n2881_));
  AND2_X1   g2689(.A1(new_n2880_), .A2(new_n2881_), .ZN(new_n2882_));
  NOR2_X1   g2690(.A1(new_n1657_), .A2(new_n1622_), .ZN(new_n2883_));
  XNOR2_X1  g2691(.A(new_n2882_), .B(new_n2883_), .ZN(new_n2884_));
  NAND2_X1  g2692(.A1(new_n2850_), .A2(new_n2860_), .ZN(new_n2885_));
  NAND2_X1  g2693(.A1(new_n2863_), .A2(new_n2885_), .ZN(new_n2886_));
  XOR2_X1   g2694(.A(new_n2884_), .B(new_n2886_), .Z(new_n2887_));
  NAND3_X1  g2695(.A1(new_n2847_), .A2(new_n2836_), .A3(new_n2871_), .ZN(new_n2888_));
  NAND2_X1  g2696(.A1(new_n2888_), .A2(new_n2870_), .ZN(new_n2889_));
  NAND2_X1  g2697(.A1(new_n2835_), .A2(new_n2870_), .ZN(new_n2890_));
  INV_X1    g2698(.A(new_n2837_), .ZN(new_n2891_));
  AOI21_X1  g2699(.A(new_n2890_), .B1(new_n2844_), .B2(new_n2891_), .ZN(new_n2892_));
  NAND2_X1  g2700(.A1(new_n2887_), .A2(new_n2869_), .ZN(new_n2893_));
  OAI22_X1  g2701(.A1(new_n2887_), .A2(new_n2889_), .B1(new_n2892_), .B2(new_n2893_), .ZN(G6280gat));
  NAND2_X1  g2702(.A1(new_n2884_), .A2(new_n2886_), .ZN(new_n2895_));
  OAI21_X1  g2703(.A(new_n2895_), .B1(new_n2892_), .B2(new_n2893_), .ZN(new_n2896_));
  OAI21_X1  g2704(.A(new_n2881_), .B1(new_n2879_), .B2(new_n2883_), .ZN(new_n2897_));
  OR2_X1    g2705(.A1(new_n2897_), .A2(KEYINPUT127), .ZN(new_n2898_));
  NOR2_X1   g2706(.A1(new_n1823_), .A2(new_n1622_), .ZN(new_n2899_));
  NAND2_X1  g2707(.A1(new_n2897_), .A2(KEYINPUT127), .ZN(new_n2900_));
  AND3_X1   g2708(.A1(new_n2898_), .A2(new_n2899_), .A3(new_n2900_), .ZN(new_n2901_));
  AOI21_X1  g2709(.A(new_n2899_), .B1(new_n2898_), .B2(new_n2900_), .ZN(new_n2902_));
  NOR2_X1   g2710(.A1(new_n2901_), .A2(new_n2902_), .ZN(new_n2903_));
  INV_X1    g2711(.A(new_n2903_), .ZN(new_n2904_));
  INV_X1    g2712(.A(new_n2899_), .ZN(new_n2905_));
  AOI22_X1  g2713(.A1(new_n2896_), .A2(new_n2904_), .B1(new_n2905_), .B2(new_n2897_), .ZN(G6287gat));
  NAND2_X1  g2714(.A1(new_n2889_), .A2(new_n2887_), .ZN(new_n2907_));
  AOI21_X1  g2715(.A(new_n2903_), .B1(new_n2886_), .B2(new_n2884_), .ZN(new_n2908_));
  AOI22_X1  g2716(.A1(new_n2896_), .A2(new_n2903_), .B1(new_n2907_), .B2(new_n2908_), .ZN(G6288gat));
endmodule


