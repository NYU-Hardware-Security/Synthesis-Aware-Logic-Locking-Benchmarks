//Secret key is'1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_c3540" written by ABC on Sun Nov 20 19:50:25 2022

module locked_c3540 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G13, G20, G33, G41, G45, G50, G58, G68,
    G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150,
    G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244,
    G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326,
    G329, G330, G343, G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G13, G20, G33, G41, G45,
    G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201_, new_n202_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1238_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201_));
  INV_X1    g0001(.A(G77), .ZN(new_n202_));
  AND2_X1   g0002(.A1(new_n201_), .A2(new_n202_), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0004(.A(G50), .B1(G58), .B2(G68), .ZN(new_n205_));
  XOR2_X1   g0005(.A(new_n205_), .B(KEYINPUT3), .Z(new_n206_));
  AND2_X1   g0006(.A1(G1), .A2(G13), .ZN(new_n207_));
  NAND3_X1  g0007(.A1(new_n206_), .A2(G20), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209_));
  NOR2_X1   g0009(.A1(new_n209_), .A2(G13), .ZN(new_n210_));
  INV_X1    g0010(.A(new_n210_), .ZN(new_n211_));
  OAI21_X1  g0011(.A(G250), .B1(G257), .B2(G264), .ZN(new_n212_));
  OAI21_X1  g0012(.A(new_n208_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g0013(.A(G107), .ZN(new_n214_));
  INV_X1    g0014(.A(G264), .ZN(new_n215_));
  NOR2_X1   g0015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g0016(.A(G68), .ZN(new_n217_));
  INV_X1    g0017(.A(G238), .ZN(new_n218_));
  INV_X1    g0018(.A(G87), .ZN(new_n219_));
  INV_X1    g0019(.A(G250), .ZN(new_n220_));
  OAI22_X1  g0020(.A1(new_n217_), .A2(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AOI211_X1 g0021(.A(new_n216_), .B(new_n221_), .C1(G116), .C2(G270), .ZN(new_n222_));
  XNOR2_X1  g0022(.A(KEYINPUT1), .B(G97), .ZN(new_n223_));
  INV_X1    g0023(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g0024(.A1(KEYINPUT2), .A2(G257), .ZN(new_n225_));
  AND2_X1   g0025(.A1(KEYINPUT2), .A2(G257), .ZN(new_n226_));
  OR3_X1    g0026(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n228_));
  INV_X1    g0028(.A(G226), .ZN(new_n229_));
  NAND2_X1  g0029(.A1(new_n229_), .A2(KEYINPUT0), .ZN(new_n230_));
  INV_X1    g0030(.A(KEYINPUT0), .ZN(new_n231_));
  NAND2_X1  g0031(.A1(new_n231_), .A2(G226), .ZN(new_n232_));
  NAND3_X1  g0032(.A1(new_n230_), .A2(new_n232_), .A3(G50), .ZN(new_n233_));
  NAND4_X1  g0033(.A1(new_n222_), .A2(new_n227_), .A3(new_n228_), .A4(new_n233_), .ZN(new_n234_));
  AOI21_X1  g0034(.A(new_n213_), .B1(new_n234_), .B2(new_n209_), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236_));
  XNOR2_X1  g0036(.A(KEYINPUT4), .B(KEYINPUT5), .ZN(new_n237_));
  XNOR2_X1  g0037(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239_));
  XNOR2_X1  g0039(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241_));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242_));
  XNOR2_X1  g0042(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XOR2_X1   g0043(.A(new_n240_), .B(new_n243_), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245_));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246_));
  XNOR2_X1  g0046(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248_));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249_));
  XNOR2_X1  g0049(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XOR2_X1   g0050(.A(new_n247_), .B(new_n250_), .Z(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252_));
  NAND3_X1  g0052(.A1(new_n252_), .A2(G13), .A3(G20), .ZN(new_n253_));
  INV_X1    g0053(.A(KEYINPUT9), .ZN(new_n254_));
  NAND2_X1  g0054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g0055(.A1(new_n252_), .A2(KEYINPUT9), .A3(G13), .A4(G20), .ZN(new_n256_));
  NAND2_X1  g0056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g0057(.A1(G1), .A2(G13), .ZN(new_n258_));
  NAND2_X1  g0058(.A1(new_n258_), .A2(KEYINPUT10), .ZN(new_n259_));
  INV_X1    g0059(.A(KEYINPUT10), .ZN(new_n260_));
  NAND3_X1  g0060(.A1(new_n260_), .A2(G1), .A3(G13), .ZN(new_n261_));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262_));
  AND3_X1   g0062(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g0063(.A1(new_n257_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g0064(.A(G58), .ZN(new_n265_));
  INV_X1    g0065(.A(G20), .ZN(new_n266_));
  NOR2_X1   g0066(.A1(new_n266_), .A2(G1), .ZN(new_n267_));
  NOR3_X1   g0067(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g0068(.A1(new_n266_), .A2(G33), .A3(G68), .ZN(new_n269_));
  INV_X1    g0069(.A(KEYINPUT28), .ZN(new_n270_));
  XNOR2_X1  g0070(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g0071(.A(G58), .B(G68), .ZN(new_n272_));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273_));
  AOI22_X1  g0073(.A1(new_n272_), .A2(G20), .B1(G159), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g0074(.A(new_n263_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g0075(.A(KEYINPUT29), .B1(new_n268_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g0076(.A1(new_n271_), .A2(new_n274_), .ZN(new_n277_));
  NAND3_X1  g0077(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n278_));
  NAND2_X1  g0078(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g0079(.A(new_n278_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n280_));
  INV_X1    g0080(.A(new_n267_), .ZN(new_n281_));
  NAND3_X1  g0081(.A1(new_n280_), .A2(G58), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g0082(.A(KEYINPUT29), .ZN(new_n283_));
  NAND3_X1  g0083(.A1(new_n279_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  AND2_X1   g0084(.A1(new_n255_), .A2(new_n256_), .ZN(new_n285_));
  AOI22_X1  g0085(.A1(new_n276_), .A2(new_n284_), .B1(new_n265_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g0086(.A(new_n252_), .B1(G41), .B2(G45), .ZN(new_n287_));
  INV_X1    g0087(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g0088(.A(KEYINPUT8), .ZN(new_n289_));
  AND2_X1   g0089(.A1(G33), .A2(G41), .ZN(new_n290_));
  OAI21_X1  g0090(.A(new_n289_), .B1(new_n290_), .B2(new_n258_), .ZN(new_n291_));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292_));
  NAND3_X1  g0092(.A1(new_n207_), .A2(KEYINPUT8), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g0093(.A(new_n288_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g0094(.A1(new_n294_), .A2(G232), .ZN(new_n295_));
  NOR2_X1   g0095(.A1(G33), .A2(G1698), .ZN(new_n296_));
  AOI22_X1  g0096(.A1(new_n296_), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n297_));
  NAND2_X1  g0097(.A1(new_n230_), .A2(new_n232_), .ZN(new_n298_));
  INV_X1    g0098(.A(G33), .ZN(new_n299_));
  NAND2_X1  g0099(.A1(new_n299_), .A2(G1698), .ZN(new_n300_));
  OAI21_X1  g0100(.A(new_n297_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g0101(.A1(new_n290_), .A2(new_n258_), .ZN(new_n302_));
  NAND2_X1  g0102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g0103(.A(G274), .ZN(new_n304_));
  NOR2_X1   g0104(.A1(new_n287_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g0105(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g0106(.A1(new_n295_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g0107(.A(G190), .ZN(new_n308_));
  NOR2_X1   g0108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g0109(.A(new_n309_), .B1(G200), .B2(new_n307_), .ZN(new_n310_));
  NAND2_X1  g0110(.A1(new_n286_), .A2(new_n310_), .ZN(new_n311_));
  OR2_X1    g0111(.A1(new_n311_), .A2(KEYINPUT30), .ZN(new_n312_));
  NOR3_X1   g0112(.A1(new_n268_), .A2(KEYINPUT29), .A3(new_n275_), .ZN(new_n313_));
  AOI21_X1  g0113(.A(new_n283_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n314_));
  OAI22_X1  g0114(.A1(new_n313_), .A2(new_n314_), .B1(G58), .B2(new_n257_), .ZN(new_n315_));
  INV_X1    g0115(.A(G179), .ZN(new_n316_));
  OR2_X1    g0116(.A1(new_n307_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g0117(.A1(new_n307_), .A2(G169), .ZN(new_n318_));
  OAI21_X1  g0118(.A(new_n317_), .B1(KEYINPUT31), .B2(new_n318_), .ZN(new_n319_));
  AND2_X1   g0119(.A1(new_n318_), .A2(KEYINPUT31), .ZN(new_n320_));
  OAI21_X1  g0120(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g0121(.A1(new_n321_), .A2(KEYINPUT30), .A3(new_n311_), .ZN(new_n322_));
  AND2_X1   g0122(.A1(new_n312_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g0123(.A(KEYINPUT27), .ZN(new_n324_));
  NOR2_X1   g0124(.A1(new_n299_), .A2(G20), .ZN(new_n325_));
  AOI22_X1  g0125(.A1(new_n325_), .A2(G58), .B1(new_n273_), .B2(G150), .ZN(new_n326_));
  OAI21_X1  g0126(.A(new_n326_), .B1(new_n266_), .B2(new_n201_), .ZN(new_n327_));
  INV_X1    g0127(.A(G50), .ZN(new_n328_));
  AOI22_X1  g0128(.A1(new_n327_), .A2(new_n278_), .B1(new_n285_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g0129(.A1(new_n280_), .A2(G50), .A3(new_n281_), .ZN(new_n330_));
  NAND2_X1  g0130(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g0131(.A1(new_n296_), .A2(G222), .ZN(new_n332_));
  INV_X1    g0132(.A(G223), .ZN(new_n333_));
  OAI221_X1 g0133(.A(new_n332_), .B1(new_n299_), .B2(new_n202_), .C1(new_n333_), .C2(new_n300_), .ZN(new_n334_));
  AOI21_X1  g0134(.A(new_n305_), .B1(new_n334_), .B2(new_n302_), .ZN(new_n335_));
  NAND2_X1  g0135(.A1(new_n294_), .A2(G226), .ZN(new_n336_));
  NAND2_X1  g0136(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g0137(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g0138(.A(new_n331_), .B1(new_n338_), .B2(G190), .ZN(new_n339_));
  NAND2_X1  g0139(.A1(new_n337_), .A2(G200), .ZN(new_n340_));
  NAND2_X1  g0140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g0141(.A(new_n341_), .B(KEYINPUT14), .ZN(new_n342_));
  INV_X1    g0142(.A(G169), .ZN(new_n343_));
  NAND2_X1  g0143(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g0144(.A(new_n344_), .B(new_n331_), .C1(G179), .C2(new_n337_), .ZN(new_n345_));
  NAND2_X1  g0145(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g0146(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g0147(.A(KEYINPUT19), .ZN(new_n348_));
  INV_X1    g0148(.A(G97), .ZN(new_n349_));
  OAI21_X1  g0149(.A(KEYINPUT17), .B1(new_n299_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351_));
  NAND3_X1  g0151(.A1(new_n351_), .A2(G33), .A3(G97), .ZN(new_n352_));
  INV_X1    g0152(.A(G232), .ZN(new_n353_));
  OAI211_X1 g0153(.A(new_n350_), .B(new_n352_), .C1(new_n353_), .C2(new_n300_), .ZN(new_n354_));
  AND3_X1   g0154(.A1(new_n230_), .A2(new_n232_), .A3(new_n296_), .ZN(new_n355_));
  OAI21_X1  g0155(.A(new_n302_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g0156(.A1(new_n291_), .A2(new_n293_), .ZN(new_n357_));
  NAND3_X1  g0157(.A1(new_n357_), .A2(G238), .A3(new_n287_), .ZN(new_n358_));
  NAND4_X1  g0158(.A1(new_n356_), .A2(new_n358_), .A3(G190), .A4(new_n306_), .ZN(new_n359_));
  NAND3_X1  g0159(.A1(new_n255_), .A2(new_n217_), .A3(new_n256_), .ZN(new_n360_));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361_));
  XNOR2_X1  g0161(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  AOI21_X1  g0162(.A(G20), .B1(G33), .B2(G77), .ZN(new_n363_));
  NAND2_X1  g0163(.A1(new_n299_), .A2(G50), .ZN(new_n364_));
  AOI22_X1  g0164(.A1(new_n363_), .A2(new_n364_), .B1(G20), .B2(G68), .ZN(new_n365_));
  NAND2_X1  g0165(.A1(new_n365_), .A2(new_n278_), .ZN(new_n366_));
  INV_X1    g0166(.A(KEYINPUT15), .ZN(new_n367_));
  NAND2_X1  g0167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g0168(.A1(new_n365_), .A2(new_n278_), .A3(KEYINPUT15), .ZN(new_n369_));
  NAND2_X1  g0169(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g0170(.A1(new_n280_), .A2(G68), .A3(new_n281_), .ZN(new_n371_));
  NAND4_X1  g0171(.A1(new_n359_), .A2(new_n362_), .A3(new_n370_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373_));
  NAND3_X1  g0173(.A1(new_n356_), .A2(new_n358_), .A3(new_n306_), .ZN(new_n374_));
  AOI21_X1  g0174(.A(new_n373_), .B1(new_n374_), .B2(G200), .ZN(new_n375_));
  INV_X1    g0175(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g0176(.A1(new_n374_), .A2(new_n373_), .A3(G200), .ZN(new_n377_));
  AOI21_X1  g0177(.A(new_n372_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g0178(.A1(new_n362_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n379_));
  NAND2_X1  g0179(.A1(new_n374_), .A2(new_n343_), .ZN(new_n380_));
  NAND4_X1  g0180(.A1(new_n356_), .A2(new_n358_), .A3(new_n316_), .A4(new_n306_), .ZN(new_n381_));
  NAND3_X1  g0181(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g0182(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g0183(.A(new_n348_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g0184(.A(new_n379_), .ZN(new_n385_));
  AND3_X1   g0185(.A1(new_n374_), .A2(new_n373_), .A3(G200), .ZN(new_n386_));
  OAI211_X1 g0186(.A(new_n385_), .B(new_n359_), .C1(new_n386_), .C2(new_n375_), .ZN(new_n387_));
  NAND3_X1  g0187(.A1(new_n387_), .A2(KEYINPUT19), .A3(new_n382_), .ZN(new_n388_));
  NAND2_X1  g0188(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g0189(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g0190(.A1(new_n347_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g0191(.A1(new_n285_), .A2(new_n202_), .ZN(new_n392_));
  NAND3_X1  g0192(.A1(new_n280_), .A2(G77), .A3(new_n281_), .ZN(new_n393_));
  XNOR2_X1  g0193(.A(KEYINPUT20), .B(G87), .ZN(new_n394_));
  NAND2_X1  g0194(.A1(new_n394_), .A2(new_n325_), .ZN(new_n395_));
  INV_X1    g0195(.A(KEYINPUT21), .ZN(new_n396_));
  NAND2_X1  g0196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g0197(.A1(new_n394_), .A2(KEYINPUT21), .A3(new_n325_), .ZN(new_n398_));
  AOI22_X1  g0198(.A1(new_n273_), .A2(G58), .B1(G20), .B2(G77), .ZN(new_n399_));
  NAND3_X1  g0199(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g0200(.A1(new_n400_), .A2(KEYINPUT22), .A3(new_n278_), .ZN(new_n401_));
  INV_X1    g0201(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g0202(.A(KEYINPUT22), .B1(new_n400_), .B2(new_n278_), .ZN(new_n403_));
  OAI211_X1 g0203(.A(new_n392_), .B(new_n393_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  AND2_X1   g0204(.A1(KEYINPUT11), .A2(G107), .ZN(new_n405_));
  NOR2_X1   g0205(.A1(KEYINPUT11), .A2(G107), .ZN(new_n406_));
  NOR3_X1   g0206(.A1(new_n405_), .A2(new_n406_), .A3(new_n299_), .ZN(new_n407_));
  INV_X1    g0207(.A(G1698), .ZN(new_n408_));
  NAND3_X1  g0208(.A1(new_n299_), .A2(new_n408_), .A3(G232), .ZN(new_n409_));
  NAND3_X1  g0209(.A1(new_n299_), .A2(G238), .A3(G1698), .ZN(new_n410_));
  NAND2_X1  g0210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g0211(.A(KEYINPUT23), .B1(new_n407_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g0212(.A1(KEYINPUT11), .A2(G107), .ZN(new_n413_));
  NAND2_X1  g0213(.A1(KEYINPUT11), .A2(G107), .ZN(new_n414_));
  NAND3_X1  g0214(.A1(new_n413_), .A2(G33), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g0215(.A(KEYINPUT23), .ZN(new_n416_));
  NAND4_X1  g0216(.A1(new_n415_), .A2(new_n416_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n417_));
  NAND3_X1  g0217(.A1(new_n412_), .A2(new_n302_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g0218(.A(new_n305_), .B1(new_n294_), .B2(G244), .ZN(new_n419_));
  NAND2_X1  g0219(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g0220(.A1(new_n420_), .A2(KEYINPUT24), .ZN(new_n421_));
  INV_X1    g0221(.A(KEYINPUT24), .ZN(new_n422_));
  NAND3_X1  g0222(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g0223(.A(new_n343_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g0224(.A1(new_n418_), .A2(new_n419_), .A3(G179), .ZN(new_n425_));
  INV_X1    g0225(.A(KEYINPUT25), .ZN(new_n426_));
  NAND2_X1  g0226(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g0227(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT25), .A4(G179), .ZN(new_n428_));
  NAND2_X1  g0228(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g0229(.A(new_n404_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g0230(.A(KEYINPUT26), .ZN(new_n431_));
  NAND2_X1  g0231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g0232(.A(KEYINPUT26), .B(new_n404_), .C1(new_n424_), .C2(new_n429_), .ZN(new_n433_));
  NAND2_X1  g0233(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g0234(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g0235(.A(new_n404_), .ZN(new_n436_));
  INV_X1    g0236(.A(new_n423_), .ZN(new_n437_));
  AOI21_X1  g0237(.A(new_n422_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n438_));
  OAI21_X1  g0238(.A(G200), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g0239(.A(new_n436_), .B(new_n439_), .C1(new_n308_), .C2(new_n420_), .ZN(new_n440_));
  NAND2_X1  g0240(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g0241(.A(new_n324_), .B1(new_n391_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g0242(.A1(new_n346_), .A2(new_n389_), .ZN(new_n443_));
  NAND4_X1  g0243(.A1(new_n443_), .A2(KEYINPUT27), .A3(new_n435_), .A4(new_n440_), .ZN(new_n444_));
  AOI21_X1  g0244(.A(new_n323_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g0245(.A(KEYINPUT12), .ZN(new_n446_));
  NOR2_X1   g0246(.A1(new_n299_), .A2(G1), .ZN(new_n447_));
  NOR2_X1   g0247(.A1(new_n447_), .A2(new_n349_), .ZN(new_n448_));
  AOI22_X1  g0248(.A1(new_n280_), .A2(new_n448_), .B1(new_n224_), .B2(new_n285_), .ZN(new_n449_));
  OAI21_X1  g0249(.A(G97), .B1(new_n405_), .B2(new_n406_), .ZN(new_n450_));
  OAI211_X1 g0250(.A(new_n450_), .B(G20), .C1(new_n214_), .C2(new_n223_), .ZN(new_n451_));
  AOI22_X1  g0251(.A1(new_n325_), .A2(G107), .B1(new_n273_), .B2(G77), .ZN(new_n452_));
  AOI21_X1  g0252(.A(new_n263_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g0253(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g0254(.A(G41), .ZN(new_n455_));
  NAND3_X1  g0255(.A1(new_n252_), .A2(new_n455_), .A3(G45), .ZN(new_n456_));
  INV_X1    g0256(.A(KEYINPUT7), .ZN(new_n457_));
  NAND2_X1  g0257(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g0258(.A(G45), .ZN(new_n459_));
  NOR3_X1   g0259(.A1(new_n459_), .A2(G1), .A3(G41), .ZN(new_n460_));
  NAND2_X1  g0260(.A1(new_n460_), .A2(KEYINPUT7), .ZN(new_n461_));
  NAND4_X1  g0261(.A1(new_n357_), .A2(G274), .A3(new_n458_), .A4(new_n461_), .ZN(new_n462_));
  NAND3_X1  g0262(.A1(new_n299_), .A2(new_n408_), .A3(G244), .ZN(new_n463_));
  NAND3_X1  g0263(.A1(new_n299_), .A2(G250), .A3(G1698), .ZN(new_n464_));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465_));
  NAND3_X1  g0265(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g0266(.A1(new_n466_), .A2(new_n302_), .ZN(new_n467_));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468_));
  NAND2_X1  g0268(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g0269(.A1(new_n290_), .A2(new_n289_), .A3(new_n258_), .ZN(new_n470_));
  AOI21_X1  g0270(.A(KEYINPUT8), .B1(new_n207_), .B2(new_n292_), .ZN(new_n471_));
  OAI211_X1 g0271(.A(G257), .B(new_n456_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g0272(.A1(new_n466_), .A2(KEYINPUT6), .A3(new_n302_), .ZN(new_n473_));
  NAND4_X1  g0273(.A1(new_n462_), .A2(new_n469_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  OAI211_X1 g0274(.A(new_n449_), .B(new_n454_), .C1(new_n474_), .C2(new_n308_), .ZN(new_n475_));
  INV_X1    g0275(.A(G200), .ZN(new_n476_));
  INV_X1    g0276(.A(new_n473_), .ZN(new_n477_));
  AOI21_X1  g0277(.A(KEYINPUT6), .B1(new_n466_), .B2(new_n302_), .ZN(new_n478_));
  NOR2_X1   g0278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AND2_X1   g0279(.A1(new_n461_), .A2(new_n458_), .ZN(new_n480_));
  AOI21_X1  g0280(.A(new_n304_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n481_));
  AOI21_X1  g0281(.A(new_n460_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n482_));
  AOI22_X1  g0282(.A1(new_n480_), .A2(new_n481_), .B1(new_n482_), .B2(G257), .ZN(new_n483_));
  AOI21_X1  g0283(.A(new_n476_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g0284(.A(new_n446_), .B1(new_n475_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g0285(.A1(new_n474_), .A2(G200), .ZN(new_n486_));
  NAND3_X1  g0286(.A1(new_n479_), .A2(new_n483_), .A3(G190), .ZN(new_n487_));
  INV_X1    g0287(.A(new_n448_), .ZN(new_n488_));
  OAI22_X1  g0288(.A1(new_n264_), .A2(new_n488_), .B1(new_n223_), .B2(new_n257_), .ZN(new_n489_));
  NOR2_X1   g0289(.A1(new_n489_), .A2(new_n453_), .ZN(new_n490_));
  NAND4_X1  g0290(.A1(new_n486_), .A2(new_n487_), .A3(new_n490_), .A4(KEYINPUT12), .ZN(new_n491_));
  INV_X1    g0291(.A(KEYINPUT13), .ZN(new_n492_));
  NAND2_X1  g0292(.A1(new_n451_), .A2(new_n452_), .ZN(new_n493_));
  AOI21_X1  g0293(.A(new_n492_), .B1(new_n493_), .B2(new_n278_), .ZN(new_n494_));
  AOI211_X1 g0294(.A(KEYINPUT13), .B(new_n263_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n495_));
  OAI21_X1  g0295(.A(new_n449_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g0296(.A1(new_n474_), .A2(new_n343_), .ZN(new_n497_));
  NAND3_X1  g0297(.A1(new_n479_), .A2(new_n483_), .A3(new_n316_), .ZN(new_n498_));
  AND2_X1   g0298(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI22_X1  g0299(.A1(new_n485_), .A2(new_n491_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g0300(.A(new_n447_), .ZN(new_n501_));
  NAND3_X1  g0301(.A1(new_n280_), .A2(new_n394_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g0302(.A(KEYINPUT35), .ZN(new_n503_));
  AOI21_X1  g0303(.A(G20), .B1(G33), .B2(G97), .ZN(new_n504_));
  OAI21_X1  g0304(.A(new_n504_), .B1(G33), .B2(new_n217_), .ZN(new_n505_));
  NAND3_X1  g0305(.A1(new_n219_), .A2(new_n349_), .A3(new_n214_), .ZN(new_n506_));
  OAI211_X1 g0306(.A(new_n278_), .B(new_n505_), .C1(new_n266_), .C2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g0307(.A1(new_n502_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g0308(.A(new_n394_), .ZN(new_n509_));
  NAND2_X1  g0309(.A1(new_n285_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g0310(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g0311(.A(new_n503_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n512_));
  OR2_X1    g0312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g0313(.A1(new_n459_), .A2(G1), .ZN(new_n514_));
  NOR2_X1   g0314(.A1(new_n514_), .A2(new_n220_), .ZN(new_n515_));
  NAND3_X1  g0315(.A1(new_n299_), .A2(G244), .A3(G1698), .ZN(new_n516_));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517_));
  NAND2_X1  g0317(.A1(new_n299_), .A2(new_n408_), .ZN(new_n518_));
  OAI211_X1 g0318(.A(new_n516_), .B(new_n517_), .C1(new_n518_), .C2(new_n218_), .ZN(new_n519_));
  AOI22_X1  g0319(.A1(new_n357_), .A2(new_n515_), .B1(new_n519_), .B2(new_n302_), .ZN(new_n520_));
  OAI211_X1 g0320(.A(G274), .B(new_n514_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n521_));
  INV_X1    g0321(.A(KEYINPUT32), .ZN(new_n522_));
  NOR2_X1   g0322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g0323(.A(KEYINPUT32), .B1(new_n481_), .B2(new_n514_), .ZN(new_n524_));
  OAI21_X1  g0324(.A(new_n520_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g0325(.A(KEYINPUT33), .ZN(new_n526_));
  NAND2_X1  g0326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g0327(.A(new_n515_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n528_));
  NAND2_X1  g0328(.A1(new_n519_), .A2(new_n302_), .ZN(new_n529_));
  NAND2_X1  g0329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g0330(.A1(new_n521_), .A2(new_n522_), .ZN(new_n531_));
  NAND3_X1  g0331(.A1(new_n481_), .A2(KEYINPUT32), .A3(new_n514_), .ZN(new_n532_));
  AOI21_X1  g0332(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g0333(.A1(new_n533_), .A2(KEYINPUT33), .ZN(new_n534_));
  AOI21_X1  g0334(.A(new_n343_), .B1(new_n527_), .B2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g0335(.A(G179), .B(new_n520_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n536_));
  INV_X1    g0336(.A(KEYINPUT34), .ZN(new_n537_));
  NAND2_X1  g0337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g0338(.A1(new_n533_), .A2(KEYINPUT34), .A3(G179), .ZN(new_n539_));
  NAND2_X1  g0339(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g0340(.A(new_n513_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  AOI211_X1 g0341(.A(new_n526_), .B(new_n530_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n542_));
  NAND2_X1  g0342(.A1(new_n531_), .A2(new_n532_), .ZN(new_n543_));
  AOI21_X1  g0343(.A(KEYINPUT33), .B1(new_n543_), .B2(new_n520_), .ZN(new_n544_));
  OAI21_X1  g0344(.A(G200), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g0345(.A1(new_n280_), .A2(G87), .A3(new_n501_), .ZN(new_n546_));
  NAND3_X1  g0346(.A1(new_n546_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n547_));
  AOI21_X1  g0347(.A(new_n547_), .B1(G190), .B2(new_n533_), .ZN(new_n548_));
  NAND2_X1  g0348(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g0349(.A1(new_n500_), .A2(new_n541_), .A3(new_n549_), .ZN(new_n550_));
  NAND3_X1  g0350(.A1(new_n299_), .A2(new_n408_), .A3(G250), .ZN(new_n551_));
  NAND3_X1  g0351(.A1(new_n299_), .A2(G257), .A3(G1698), .ZN(new_n552_));
  NAND2_X1  g0352(.A1(G33), .A2(G294), .ZN(new_n553_));
  NAND3_X1  g0353(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g0354(.A(KEYINPUT40), .ZN(new_n555_));
  AND3_X1   g0355(.A1(new_n554_), .A2(new_n555_), .A3(new_n302_), .ZN(new_n556_));
  AOI21_X1  g0356(.A(new_n555_), .B1(new_n554_), .B2(new_n302_), .ZN(new_n557_));
  OAI21_X1  g0357(.A(new_n462_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g0358(.A1(new_n482_), .A2(G264), .ZN(new_n559_));
  NAND2_X1  g0359(.A1(new_n559_), .A2(G179), .ZN(new_n560_));
  OAI21_X1  g0360(.A(KEYINPUT41), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g0361(.A(new_n559_), .B(new_n462_), .C1(new_n557_), .C2(new_n556_), .ZN(new_n562_));
  NAND2_X1  g0362(.A1(new_n562_), .A2(G169), .ZN(new_n563_));
  INV_X1    g0363(.A(new_n557_), .ZN(new_n564_));
  NAND3_X1  g0364(.A1(new_n554_), .A2(new_n555_), .A3(new_n302_), .ZN(new_n565_));
  NAND2_X1  g0365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g0366(.A(KEYINPUT41), .ZN(new_n567_));
  AOI21_X1  g0367(.A(new_n316_), .B1(new_n482_), .B2(G264), .ZN(new_n568_));
  NAND4_X1  g0368(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .A4(new_n462_), .ZN(new_n569_));
  NAND3_X1  g0369(.A1(new_n561_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g0370(.A1(new_n299_), .A2(G87), .ZN(new_n571_));
  AOI21_X1  g0371(.A(G20), .B1(new_n571_), .B2(new_n517_), .ZN(new_n572_));
  NAND2_X1  g0372(.A1(new_n278_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g0373(.A1(new_n501_), .A2(G107), .ZN(new_n574_));
  OAI21_X1  g0374(.A(new_n573_), .B1(new_n264_), .B2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g0375(.A1(new_n405_), .A2(new_n406_), .ZN(new_n576_));
  INV_X1    g0376(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g0377(.A(new_n577_), .B1(KEYINPUT9), .B2(G20), .ZN(new_n578_));
  NOR2_X1   g0378(.A1(new_n280_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g0379(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g0380(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g0381(.A1(new_n570_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g0382(.A(KEYINPUT42), .ZN(new_n583_));
  NAND2_X1  g0383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g0384(.A1(new_n570_), .A2(KEYINPUT42), .A3(new_n581_), .ZN(new_n585_));
  OR2_X1    g0385(.A1(new_n562_), .A2(new_n308_), .ZN(new_n586_));
  NAND2_X1  g0386(.A1(new_n562_), .A2(G200), .ZN(new_n587_));
  NAND3_X1  g0387(.A1(new_n586_), .A2(new_n580_), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g0388(.A1(new_n584_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  NOR2_X1   g0389(.A1(new_n550_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g0390(.A1(new_n357_), .A2(G270), .A3(new_n456_), .ZN(new_n591_));
  NOR3_X1   g0391(.A1(new_n518_), .A2(new_n226_), .A3(new_n225_), .ZN(new_n592_));
  INV_X1    g0392(.A(G303), .ZN(new_n593_));
  OAI22_X1  g0393(.A1(new_n300_), .A2(new_n215_), .B1(new_n299_), .B2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g0394(.A(new_n302_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g0395(.A1(new_n462_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g0396(.A1(new_n596_), .A2(G200), .ZN(new_n597_));
  XNOR2_X1  g0397(.A(new_n597_), .B(KEYINPUT39), .ZN(new_n598_));
  NAND2_X1  g0398(.A1(new_n349_), .A2(KEYINPUT1), .ZN(new_n599_));
  INV_X1    g0399(.A(KEYINPUT1), .ZN(new_n600_));
  NAND2_X1  g0400(.A1(new_n600_), .A2(G97), .ZN(new_n601_));
  NAND3_X1  g0401(.A1(new_n599_), .A2(new_n601_), .A3(new_n273_), .ZN(new_n602_));
  NAND3_X1  g0402(.A1(new_n266_), .A2(G33), .A3(G283), .ZN(new_n603_));
  INV_X1    g0403(.A(KEYINPUT36), .ZN(new_n604_));
  NAND2_X1  g0404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g0405(.A1(G20), .A2(G116), .ZN(new_n606_));
  NAND4_X1  g0406(.A1(new_n266_), .A2(KEYINPUT36), .A3(G33), .A4(G283), .ZN(new_n607_));
  NAND4_X1  g0407(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g0408(.A1(new_n608_), .A2(new_n278_), .ZN(new_n609_));
  NAND4_X1  g0409(.A1(new_n257_), .A2(new_n263_), .A3(G116), .A4(new_n501_), .ZN(new_n610_));
  INV_X1    g0410(.A(G116), .ZN(new_n611_));
  NAND2_X1  g0411(.A1(new_n285_), .A2(new_n611_), .ZN(new_n612_));
  AND3_X1   g0412(.A1(new_n609_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g0413(.A(new_n613_), .B1(new_n308_), .B2(new_n596_), .ZN(new_n614_));
  NOR2_X1   g0414(.A1(new_n598_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g0415(.A1(new_n609_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n616_));
  NAND3_X1  g0416(.A1(new_n616_), .A2(new_n596_), .A3(G169), .ZN(new_n617_));
  NAND4_X1  g0417(.A1(new_n462_), .A2(new_n591_), .A3(G179), .A4(new_n595_), .ZN(new_n618_));
  INV_X1    g0418(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g0419(.A(KEYINPUT37), .B1(new_n619_), .B2(new_n616_), .ZN(new_n620_));
  INV_X1    g0420(.A(KEYINPUT37), .ZN(new_n621_));
  NOR3_X1   g0421(.A1(new_n613_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g0422(.A(new_n617_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g0423(.A(KEYINPUT38), .ZN(new_n624_));
  NAND2_X1  g0424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g0425(.A(KEYINPUT38), .B(new_n617_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n626_));
  AOI21_X1  g0426(.A(new_n615_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AND3_X1   g0427(.A1(new_n445_), .A2(new_n590_), .A3(new_n627_), .ZN(G372));
  AND3_X1   g0428(.A1(new_n500_), .A2(new_n541_), .A3(new_n549_), .ZN(new_n629_));
  AND3_X1   g0429(.A1(new_n570_), .A2(KEYINPUT42), .A3(new_n581_), .ZN(new_n630_));
  AOI21_X1  g0430(.A(KEYINPUT42), .B1(new_n570_), .B2(new_n581_), .ZN(new_n631_));
  INV_X1    g0431(.A(new_n588_), .ZN(new_n632_));
  NOR3_X1   g0432(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND3_X1  g0433(.A1(new_n629_), .A2(new_n633_), .A3(new_n623_), .ZN(new_n634_));
  NAND2_X1  g0434(.A1(new_n584_), .A2(new_n585_), .ZN(new_n635_));
  NAND2_X1  g0435(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g0436(.A1(new_n511_), .A2(new_n512_), .ZN(new_n637_));
  AND2_X1   g0437(.A1(new_n538_), .A2(new_n539_), .ZN(new_n638_));
  OAI21_X1  g0438(.A(G169), .B1(new_n542_), .B2(new_n544_), .ZN(new_n639_));
  AOI21_X1  g0439(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g0440(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n641_));
  AOI21_X1  g0441(.A(new_n641_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n642_));
  NOR2_X1   g0442(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g0443(.A1(new_n634_), .A2(new_n636_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g0444(.A1(new_n445_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g0445(.A(new_n382_), .B(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g0446(.A(new_n646_), .B1(new_n390_), .B2(new_n434_), .ZN(new_n647_));
  OAI21_X1  g0447(.A(new_n321_), .B1(new_n647_), .B2(new_n323_), .ZN(new_n648_));
  NAND2_X1  g0448(.A1(new_n648_), .A2(new_n342_), .ZN(new_n649_));
  AND2_X1   g0449(.A1(new_n649_), .A2(new_n345_), .ZN(new_n650_));
  NAND2_X1  g0450(.A1(new_n645_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g0451(.A(new_n651_), .B(KEYINPUT44), .Z(G369));
  INV_X1    g0452(.A(G13), .ZN(new_n653_));
  INV_X1    g0453(.A(G213), .ZN(new_n654_));
  NOR4_X1   g0454(.A1(new_n653_), .A2(new_n654_), .A3(G1), .A4(G20), .ZN(new_n655_));
  INV_X1    g0455(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g0456(.A(G343), .ZN(new_n657_));
  NOR2_X1   g0457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g0458(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g0459(.A1(new_n580_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g0460(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g0461(.A1(new_n633_), .A2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g0462(.A(KEYINPUT45), .B(KEYINPUT46), .Z(new_n663_));
  INV_X1    g0463(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g0464(.A1(new_n635_), .A2(new_n660_), .ZN(new_n665_));
  AND3_X1   g0465(.A1(new_n662_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g0466(.A(new_n664_), .B1(new_n662_), .B2(new_n665_), .ZN(new_n667_));
  OR2_X1    g0467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g0468(.A1(new_n625_), .A2(new_n626_), .ZN(new_n669_));
  NOR2_X1   g0469(.A1(new_n613_), .A2(new_n659_), .ZN(new_n670_));
  MUX2_X1   g0470(.A(new_n627_), .B(new_n669_), .S(new_n670_), .Z(new_n671_));
  XNOR2_X1  g0471(.A(KEYINPUT47), .B(G330), .ZN(new_n672_));
  NAND3_X1  g0472(.A1(new_n668_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g0473(.A(new_n669_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n674_));
  NOR2_X1   g0474(.A1(new_n630_), .A2(new_n631_), .ZN(new_n675_));
  AND2_X1   g0475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g0476(.A(new_n673_), .B1(new_n676_), .B2(new_n658_), .ZN(G399));
  INV_X1    g0477(.A(KEYINPUT48), .ZN(new_n678_));
  OAI21_X1  g0478(.A(new_n678_), .B1(new_n211_), .B2(G41), .ZN(new_n679_));
  NAND3_X1  g0479(.A1(new_n210_), .A2(KEYINPUT48), .A3(new_n455_), .ZN(new_n680_));
  NAND2_X1  g0480(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NOR3_X1   g0481(.A1(new_n681_), .A2(KEYINPUT49), .A3(new_n252_), .ZN(new_n682_));
  NOR2_X1   g0482(.A1(new_n506_), .A2(G116), .ZN(new_n683_));
  INV_X1    g0483(.A(new_n683_), .ZN(new_n684_));
  NOR2_X1   g0484(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g0485(.A(KEYINPUT49), .B1(new_n681_), .B2(new_n252_), .ZN(new_n686_));
  AOI22_X1  g0486(.A1(new_n685_), .A2(new_n686_), .B1(new_n206_), .B2(new_n681_), .ZN(new_n687_));
  NAND4_X1  g0487(.A1(new_n629_), .A2(new_n633_), .A3(new_n627_), .A4(new_n659_), .ZN(new_n688_));
  INV_X1    g0488(.A(KEYINPUT51), .ZN(new_n689_));
  AND3_X1   g0489(.A1(new_n474_), .A2(new_n316_), .A3(new_n596_), .ZN(new_n690_));
  OAI211_X1 g0490(.A(new_n562_), .B(new_n690_), .C1(new_n542_), .C2(new_n544_), .ZN(new_n691_));
  NOR3_X1   g0491(.A1(new_n562_), .A2(new_n474_), .A3(new_n618_), .ZN(new_n692_));
  NAND3_X1  g0492(.A1(new_n692_), .A2(new_n527_), .A3(new_n534_), .ZN(new_n693_));
  NAND2_X1  g0493(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g0494(.A(new_n689_), .B1(new_n694_), .B2(new_n658_), .ZN(new_n695_));
  NAND2_X1  g0495(.A1(new_n688_), .A2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g0496(.A1(new_n590_), .A2(new_n689_), .A3(new_n627_), .A4(new_n659_), .ZN(new_n697_));
  AND2_X1   g0497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g0498(.A1(new_n698_), .A2(G330), .ZN(new_n699_));
  INV_X1    g0499(.A(new_n623_), .ZN(new_n700_));
  NOR3_X1   g0500(.A1(new_n550_), .A2(new_n589_), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g0501(.A(new_n643_), .B1(new_n550_), .B2(new_n675_), .ZN(new_n702_));
  OAI21_X1  g0502(.A(new_n659_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g0503(.A(KEYINPUT50), .ZN(new_n704_));
  NAND2_X1  g0504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g0505(.A(KEYINPUT50), .B(new_n659_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g0506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g0507(.A1(new_n699_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g0508(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g0509(.A(new_n687_), .B1(new_n709_), .B2(G1), .ZN(G364));
  XNOR2_X1  g0510(.A(new_n671_), .B(G330), .ZN(new_n711_));
  XNOR2_X1  g0511(.A(new_n711_), .B(KEYINPUT52), .ZN(new_n712_));
  NAND2_X1  g0512(.A1(new_n712_), .A2(new_n681_), .ZN(new_n713_));
  XOR2_X1   g0513(.A(new_n713_), .B(KEYINPUT53), .Z(new_n714_));
  NOR2_X1   g0514(.A1(new_n653_), .A2(G20), .ZN(new_n715_));
  AOI21_X1  g0515(.A(new_n252_), .B1(new_n715_), .B2(G45), .ZN(new_n716_));
  XNOR2_X1  g0516(.A(new_n716_), .B(KEYINPUT54), .ZN(new_n717_));
  INV_X1    g0517(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g0518(.A1(new_n712_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g0519(.A1(new_n718_), .A2(new_n681_), .ZN(new_n720_));
  INV_X1    g0520(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g0521(.A(new_n258_), .B1(G20), .B2(new_n343_), .ZN(new_n722_));
  OR2_X1    g0522(.A1(new_n722_), .A2(KEYINPUT60), .ZN(new_n723_));
  NAND2_X1  g0523(.A1(new_n722_), .A2(KEYINPUT60), .ZN(new_n724_));
  NAND2_X1  g0524(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g0525(.A(new_n725_), .ZN(new_n726_));
  OR2_X1    g0526(.A1(new_n476_), .A2(KEYINPUT56), .ZN(new_n727_));
  NAND2_X1  g0527(.A1(new_n476_), .A2(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g0528(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g0529(.A(new_n729_), .ZN(new_n730_));
  NOR3_X1   g0530(.A1(new_n266_), .A2(new_n316_), .A3(new_n308_), .ZN(new_n731_));
  NAND2_X1  g0531(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g0532(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g0533(.A1(new_n731_), .A2(new_n476_), .ZN(new_n734_));
  INV_X1    g0534(.A(new_n734_), .ZN(new_n735_));
  AOI22_X1  g0535(.A1(new_n733_), .A2(G50), .B1(new_n735_), .B2(G58), .ZN(new_n736_));
  NOR2_X1   g0536(.A1(new_n266_), .A2(G190), .ZN(new_n737_));
  INV_X1    g0537(.A(new_n737_), .ZN(new_n738_));
  NOR2_X1   g0538(.A1(new_n738_), .A2(new_n316_), .ZN(new_n739_));
  NAND2_X1  g0539(.A1(new_n730_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g0540(.A1(new_n739_), .A2(new_n729_), .ZN(new_n741_));
  OAI221_X1 g0541(.A(new_n736_), .B1(new_n217_), .B2(new_n740_), .C1(new_n202_), .C2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g0542(.A(new_n742_), .B(KEYINPUT57), .Z(new_n743_));
  NOR2_X1   g0543(.A1(new_n266_), .A2(G179), .ZN(new_n744_));
  NAND3_X1  g0544(.A1(new_n730_), .A2(G190), .A3(new_n744_), .ZN(new_n745_));
  NOR2_X1   g0545(.A1(new_n745_), .A2(new_n219_), .ZN(new_n746_));
  NAND3_X1  g0546(.A1(new_n730_), .A2(new_n308_), .A3(new_n744_), .ZN(new_n747_));
  NOR2_X1   g0547(.A1(new_n747_), .A2(new_n214_), .ZN(new_n748_));
  NOR3_X1   g0548(.A1(new_n746_), .A2(new_n748_), .A3(G33), .ZN(new_n749_));
  OAI21_X1  g0549(.A(G20), .B1(G179), .B2(G200), .ZN(new_n750_));
  INV_X1    g0550(.A(KEYINPUT55), .ZN(new_n751_));
  XNOR2_X1  g0551(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  NOR2_X1   g0552(.A1(new_n752_), .A2(new_n737_), .ZN(new_n753_));
  INV_X1    g0553(.A(new_n753_), .ZN(new_n754_));
  NOR2_X1   g0554(.A1(new_n754_), .A2(new_n224_), .ZN(new_n755_));
  NOR2_X1   g0555(.A1(new_n752_), .A2(new_n738_), .ZN(new_n756_));
  AOI21_X1  g0556(.A(new_n755_), .B1(G159), .B2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g0557(.A1(new_n743_), .A2(new_n749_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g0558(.A(new_n740_), .ZN(new_n759_));
  INV_X1    g0559(.A(new_n741_), .ZN(new_n760_));
  XNOR2_X1  g0560(.A(KEYINPUT58), .B(G311), .ZN(new_n761_));
  AOI22_X1  g0561(.A1(new_n759_), .A2(G317), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g0562(.A(G294), .ZN(new_n763_));
  INV_X1    g0563(.A(G322), .ZN(new_n764_));
  OAI221_X1 g0564(.A(new_n762_), .B1(new_n763_), .B2(new_n754_), .C1(new_n764_), .C2(new_n734_), .ZN(new_n765_));
  NAND2_X1  g0565(.A1(new_n756_), .A2(G329), .ZN(new_n766_));
  XOR2_X1   g0566(.A(new_n766_), .B(KEYINPUT59), .Z(new_n767_));
  AOI21_X1  g0567(.A(new_n299_), .B1(new_n733_), .B2(G326), .ZN(new_n768_));
  INV_X1    g0568(.A(G283), .ZN(new_n769_));
  OAI221_X1 g0569(.A(new_n768_), .B1(new_n769_), .B2(new_n747_), .C1(new_n593_), .C2(new_n745_), .ZN(new_n770_));
  OR3_X1    g0570(.A1(new_n765_), .A2(new_n767_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g0571(.A(new_n726_), .B1(new_n758_), .B2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773_));
  XNOR2_X1  g0573(.A(new_n773_), .B(KEYINPUT62), .ZN(new_n774_));
  INV_X1    g0574(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g0575(.A1(new_n775_), .A2(G20), .ZN(new_n776_));
  NOR2_X1   g0576(.A1(new_n776_), .A2(new_n725_), .ZN(new_n777_));
  NOR2_X1   g0577(.A1(new_n211_), .A2(new_n299_), .ZN(new_n778_));
  INV_X1    g0578(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g0579(.A(new_n779_), .B1(new_n250_), .B2(G45), .ZN(new_n780_));
  INV_X1    g0580(.A(new_n206_), .ZN(new_n781_));
  OAI21_X1  g0581(.A(new_n780_), .B1(G45), .B2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g0582(.A(new_n782_), .B(KEYINPUT61), .Z(new_n783_));
  INV_X1    g0583(.A(G355), .ZN(new_n784_));
  NAND2_X1  g0584(.A1(new_n210_), .A2(new_n299_), .ZN(new_n785_));
  OAI221_X1 g0585(.A(new_n783_), .B1(G116), .B2(new_n210_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  AOI211_X1 g0586(.A(new_n721_), .B(new_n772_), .C1(new_n777_), .C2(new_n786_), .ZN(new_n787_));
  INV_X1    g0587(.A(new_n776_), .ZN(new_n788_));
  OAI21_X1  g0588(.A(new_n787_), .B1(new_n671_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g0589(.A1(new_n714_), .A2(new_n719_), .A3(new_n789_), .ZN(G396));
  NAND2_X1  g0590(.A1(new_n698_), .A2(new_n672_), .ZN(new_n791_));
  INV_X1    g0591(.A(new_n791_), .ZN(new_n792_));
  NAND2_X1  g0592(.A1(new_n404_), .A2(new_n658_), .ZN(new_n793_));
  INV_X1    g0593(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g0594(.A(G169), .B1(new_n437_), .B2(new_n438_), .ZN(new_n795_));
  NAND3_X1  g0595(.A1(new_n795_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n796_));
  AOI21_X1  g0596(.A(KEYINPUT26), .B1(new_n796_), .B2(new_n404_), .ZN(new_n797_));
  INV_X1    g0597(.A(new_n433_), .ZN(new_n798_));
  OAI21_X1  g0598(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g0599(.A1(new_n432_), .A2(new_n440_), .A3(new_n433_), .A4(new_n793_), .ZN(new_n800_));
  NAND2_X1  g0600(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g0601(.A1(new_n801_), .A2(KEYINPUT63), .ZN(new_n802_));
  INV_X1    g0602(.A(KEYINPUT63), .ZN(new_n803_));
  AOI21_X1  g0603(.A(new_n803_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n804_));
  NOR2_X1   g0604(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g0605(.A1(new_n705_), .A2(new_n805_), .A3(new_n706_), .ZN(new_n806_));
  INV_X1    g0606(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g0607(.A(new_n805_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n808_));
  OAI21_X1  g0608(.A(new_n792_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g0609(.A1(new_n809_), .A2(KEYINPUT64), .ZN(new_n810_));
  INV_X1    g0610(.A(KEYINPUT64), .ZN(new_n811_));
  OAI211_X1 g0611(.A(new_n792_), .B(new_n811_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g0612(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g0613(.A(new_n805_), .ZN(new_n814_));
  NAND2_X1  g0614(.A1(new_n707_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g0615(.A1(new_n815_), .A2(new_n791_), .A3(new_n806_), .ZN(new_n816_));
  INV_X1    g0616(.A(KEYINPUT65), .ZN(new_n817_));
  NAND2_X1  g0617(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g0618(.A1(new_n815_), .A2(KEYINPUT65), .A3(new_n791_), .A4(new_n806_), .ZN(new_n819_));
  NAND2_X1  g0619(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g0620(.A1(new_n813_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g0621(.A(new_n801_), .ZN(new_n822_));
  NAND2_X1  g0622(.A1(new_n822_), .A2(new_n774_), .ZN(new_n823_));
  NOR2_X1   g0623(.A1(new_n725_), .A2(new_n773_), .ZN(new_n824_));
  INV_X1    g0624(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g0625(.A(new_n720_), .B1(new_n825_), .B2(G77), .ZN(new_n826_));
  OAI22_X1  g0626(.A1(new_n732_), .A2(new_n593_), .B1(new_n734_), .B2(new_n763_), .ZN(new_n827_));
  AOI211_X1 g0627(.A(new_n827_), .B(new_n755_), .C1(G116), .C2(new_n760_), .ZN(new_n828_));
  INV_X1    g0628(.A(new_n745_), .ZN(new_n829_));
  NAND2_X1  g0629(.A1(new_n829_), .A2(G107), .ZN(new_n830_));
  OAI21_X1  g0630(.A(G33), .B1(new_n740_), .B2(new_n769_), .ZN(new_n831_));
  INV_X1    g0631(.A(new_n747_), .ZN(new_n832_));
  AOI21_X1  g0632(.A(new_n831_), .B1(G87), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g0633(.A1(new_n756_), .A2(G311), .ZN(new_n834_));
  NAND4_X1  g0634(.A1(new_n828_), .A2(new_n830_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  AOI22_X1  g0635(.A1(new_n733_), .A2(G137), .B1(new_n735_), .B2(G143), .ZN(new_n836_));
  INV_X1    g0636(.A(G150), .ZN(new_n837_));
  INV_X1    g0637(.A(G159), .ZN(new_n838_));
  OAI221_X1 g0638(.A(new_n836_), .B1(new_n837_), .B2(new_n740_), .C1(new_n838_), .C2(new_n741_), .ZN(new_n839_));
  INV_X1    g0639(.A(KEYINPUT68), .ZN(new_n840_));
  INV_X1    g0640(.A(KEYINPUT67), .ZN(new_n841_));
  OAI21_X1  g0641(.A(new_n841_), .B1(new_n745_), .B2(new_n328_), .ZN(new_n842_));
  NAND3_X1  g0642(.A1(new_n829_), .A2(KEYINPUT67), .A3(G50), .ZN(new_n843_));
  AOI22_X1  g0643(.A1(new_n839_), .A2(new_n840_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI221_X1 g0644(.A(new_n844_), .B1(new_n840_), .B2(new_n839_), .C1(new_n265_), .C2(new_n754_), .ZN(new_n845_));
  XOR2_X1   g0645(.A(new_n845_), .B(KEYINPUT69), .Z(new_n846_));
  INV_X1    g0646(.A(new_n756_), .ZN(new_n847_));
  INV_X1    g0647(.A(G132), .ZN(new_n848_));
  OAI221_X1 g0648(.A(new_n299_), .B1(new_n747_), .B2(new_n217_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g0649(.A(new_n835_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g0650(.A(new_n826_), .B1(new_n850_), .B2(new_n725_), .ZN(new_n851_));
  AOI22_X1  g0651(.A1(new_n821_), .A2(new_n681_), .B1(new_n823_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g0652(.A(KEYINPUT66), .ZN(new_n853_));
  AOI21_X1  g0653(.A(new_n853_), .B1(new_n821_), .B2(new_n718_), .ZN(new_n854_));
  AOI22_X1  g0654(.A1(new_n810_), .A2(new_n812_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n855_));
  NOR3_X1   g0655(.A1(new_n855_), .A2(KEYINPUT66), .A3(new_n717_), .ZN(new_n856_));
  OAI21_X1  g0656(.A(new_n852_), .B1(new_n854_), .B2(new_n856_), .ZN(G384));
  NAND2_X1  g0657(.A1(new_n445_), .A2(new_n698_), .ZN(new_n858_));
  INV_X1    g0658(.A(KEYINPUT71), .ZN(new_n859_));
  XOR2_X1   g0659(.A(new_n655_), .B(KEYINPUT70), .Z(new_n860_));
  INV_X1    g0660(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g0661(.A(new_n859_), .B1(new_n286_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g0662(.A1(new_n315_), .A2(KEYINPUT71), .A3(new_n860_), .ZN(new_n863_));
  NAND2_X1  g0663(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g0664(.A1(new_n312_), .A2(new_n322_), .A3(new_n864_), .ZN(new_n865_));
  NAND3_X1  g0665(.A1(new_n317_), .A2(new_n318_), .A3(new_n861_), .ZN(new_n866_));
  NAND2_X1  g0666(.A1(new_n315_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g0667(.A(new_n310_), .ZN(new_n868_));
  NAND2_X1  g0668(.A1(new_n315_), .A2(KEYINPUT72), .ZN(new_n869_));
  INV_X1    g0669(.A(KEYINPUT72), .ZN(new_n870_));
  NAND2_X1  g0670(.A1(new_n286_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g0671(.A(new_n868_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g0672(.A(KEYINPUT73), .ZN(new_n873_));
  OAI21_X1  g0673(.A(new_n867_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  AOI211_X1 g0674(.A(KEYINPUT73), .B(new_n868_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n875_));
  OAI21_X1  g0675(.A(new_n865_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g0676(.A1(new_n385_), .A2(new_n659_), .ZN(new_n877_));
  NOR3_X1   g0677(.A1(new_n378_), .A2(new_n383_), .A3(new_n348_), .ZN(new_n878_));
  AOI21_X1  g0678(.A(KEYINPUT19), .B1(new_n387_), .B2(new_n382_), .ZN(new_n879_));
  OAI21_X1  g0679(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NOR3_X1   g0680(.A1(new_n378_), .A2(new_n383_), .A3(new_n877_), .ZN(new_n881_));
  INV_X1    g0681(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g0682(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g0683(.A1(new_n876_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g0684(.A1(new_n884_), .A2(new_n822_), .ZN(new_n885_));
  NAND2_X1  g0685(.A1(new_n698_), .A2(new_n885_), .ZN(new_n886_));
  MUX2_X1   g0686(.A(new_n445_), .B(new_n858_), .S(new_n886_), .Z(new_n887_));
  XOR2_X1   g0687(.A(new_n887_), .B(KEYINPUT75), .Z(new_n888_));
  NAND2_X1  g0688(.A1(new_n888_), .A2(new_n672_), .ZN(new_n889_));
  OAI211_X1 g0689(.A(new_n659_), .B(new_n801_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n890_));
  AOI21_X1  g0690(.A(new_n658_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n891_));
  INV_X1    g0691(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g0692(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g0693(.A(new_n884_), .ZN(new_n894_));
  NAND2_X1  g0694(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g0695(.A(KEYINPUT74), .ZN(new_n896_));
  NOR2_X1   g0696(.A1(new_n321_), .A2(new_n860_), .ZN(new_n897_));
  INV_X1    g0697(.A(new_n897_), .ZN(new_n898_));
  NAND3_X1  g0698(.A1(new_n895_), .A2(new_n896_), .A3(new_n898_), .ZN(new_n899_));
  NOR2_X1   g0699(.A1(new_n382_), .A2(new_n658_), .ZN(new_n900_));
  NAND2_X1  g0700(.A1(new_n876_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g0701(.A(new_n884_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n902_));
  OAI21_X1  g0702(.A(KEYINPUT74), .B1(new_n902_), .B2(new_n897_), .ZN(new_n903_));
  NAND3_X1  g0703(.A1(new_n899_), .A2(new_n901_), .A3(new_n903_), .ZN(new_n904_));
  NAND3_X1  g0704(.A1(new_n445_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n905_));
  NAND2_X1  g0705(.A1(new_n905_), .A2(new_n650_), .ZN(new_n906_));
  XNOR2_X1  g0706(.A(new_n904_), .B(new_n906_), .ZN(new_n907_));
  OR2_X1    g0707(.A1(new_n889_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g0708(.A1(new_n889_), .A2(new_n907_), .ZN(new_n909_));
  OAI211_X1 g0709(.A(new_n908_), .B(new_n909_), .C1(new_n252_), .C2(new_n715_), .ZN(new_n910_));
  OAI21_X1  g0710(.A(G77), .B1(new_n265_), .B2(new_n217_), .ZN(new_n911_));
  OAI22_X1  g0711(.A1(new_n911_), .A2(new_n205_), .B1(G50), .B2(new_n217_), .ZN(new_n912_));
  NAND3_X1  g0712(.A1(new_n912_), .A2(G1), .A3(new_n653_), .ZN(new_n913_));
  OAI21_X1  g0713(.A(new_n450_), .B1(new_n223_), .B2(new_n214_), .ZN(new_n914_));
  NAND4_X1  g0714(.A1(new_n914_), .A2(G20), .A3(G116), .A4(new_n207_), .ZN(new_n915_));
  NAND3_X1  g0715(.A1(new_n910_), .A2(new_n913_), .A3(new_n915_), .ZN(new_n916_));
  XOR2_X1   g0716(.A(new_n916_), .B(KEYINPUT76), .Z(G367));
  INV_X1    g0717(.A(KEYINPUT80), .ZN(new_n918_));
  AND2_X1   g0718(.A1(new_n671_), .A2(G330), .ZN(new_n919_));
  NAND2_X1  g0719(.A1(new_n496_), .A2(new_n658_), .ZN(new_n920_));
  XOR2_X1   g0720(.A(new_n500_), .B(new_n920_), .Z(new_n921_));
  INV_X1    g0721(.A(new_n921_), .ZN(new_n922_));
  NAND3_X1  g0722(.A1(new_n668_), .A2(new_n919_), .A3(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g0723(.A(new_n923_), .B(KEYINPUT78), .ZN(new_n924_));
  AOI21_X1  g0724(.A(new_n921_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n925_));
  INV_X1    g0725(.A(new_n641_), .ZN(new_n926_));
  OAI21_X1  g0726(.A(new_n659_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g0727(.A1(new_n640_), .A2(new_n547_), .A3(new_n658_), .ZN(new_n928_));
  NAND2_X1  g0728(.A1(new_n547_), .A2(new_n658_), .ZN(new_n929_));
  NAND3_X1  g0729(.A1(new_n541_), .A2(new_n549_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g0730(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g0731(.A1(new_n927_), .A2(new_n931_), .ZN(new_n932_));
  INV_X1    g0732(.A(KEYINPUT79), .ZN(new_n933_));
  XNOR2_X1  g0733(.A(new_n932_), .B(new_n933_), .ZN(new_n934_));
  INV_X1    g0734(.A(new_n931_), .ZN(new_n935_));
  OAI211_X1 g0735(.A(new_n659_), .B(new_n935_), .C1(new_n925_), .C2(new_n926_), .ZN(new_n936_));
  OR2_X1    g0736(.A1(new_n936_), .A2(KEYINPUT77), .ZN(new_n937_));
  NAND2_X1  g0737(.A1(new_n936_), .A2(KEYINPUT77), .ZN(new_n938_));
  AND2_X1   g0738(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  OAI211_X1 g0739(.A(new_n918_), .B(new_n924_), .C1(new_n934_), .C2(new_n939_), .ZN(new_n940_));
  INV_X1    g0740(.A(new_n924_), .ZN(new_n941_));
  AOI22_X1  g0741(.A1(new_n937_), .A2(new_n938_), .B1(new_n941_), .B2(KEYINPUT80), .ZN(new_n942_));
  XNOR2_X1  g0742(.A(new_n932_), .B(KEYINPUT79), .ZN(new_n943_));
  OAI211_X1 g0743(.A(new_n942_), .B(new_n943_), .C1(KEYINPUT80), .C2(new_n941_), .ZN(new_n944_));
  AND3_X1   g0744(.A1(new_n940_), .A2(new_n944_), .A3(new_n681_), .ZN(new_n945_));
  XNOR2_X1  g0745(.A(new_n668_), .B(new_n919_), .ZN(new_n946_));
  NAND2_X1  g0746(.A1(new_n669_), .A2(new_n659_), .ZN(new_n947_));
  XNOR2_X1  g0747(.A(new_n946_), .B(new_n947_), .ZN(new_n948_));
  OR2_X1    g0748(.A1(new_n948_), .A2(new_n708_), .ZN(new_n949_));
  INV_X1    g0749(.A(KEYINPUT84), .ZN(new_n950_));
  AOI21_X1  g0750(.A(new_n658_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n951_));
  INV_X1    g0751(.A(new_n500_), .ZN(new_n952_));
  NAND2_X1  g0752(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g0753(.A(KEYINPUT82), .ZN(new_n954_));
  XNOR2_X1  g0754(.A(new_n953_), .B(new_n954_), .ZN(new_n955_));
  OAI211_X1 g0755(.A(KEYINPUT83), .B(new_n922_), .C1(new_n676_), .C2(new_n658_), .ZN(new_n956_));
  INV_X1    g0756(.A(KEYINPUT83), .ZN(new_n957_));
  OAI21_X1  g0757(.A(new_n957_), .B1(new_n951_), .B2(new_n921_), .ZN(new_n958_));
  NAND2_X1  g0758(.A1(new_n956_), .A2(new_n958_), .ZN(new_n959_));
  XOR2_X1   g0759(.A(new_n673_), .B(KEYINPUT81), .Z(new_n960_));
  NAND3_X1  g0760(.A1(new_n955_), .A2(new_n959_), .A3(new_n960_), .ZN(new_n961_));
  INV_X1    g0761(.A(new_n961_), .ZN(new_n962_));
  AOI21_X1  g0762(.A(new_n960_), .B1(new_n955_), .B2(new_n959_), .ZN(new_n963_));
  OAI21_X1  g0763(.A(new_n950_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  INV_X1    g0764(.A(new_n963_), .ZN(new_n965_));
  NAND3_X1  g0765(.A1(new_n965_), .A2(KEYINPUT84), .A3(new_n961_), .ZN(new_n966_));
  AOI21_X1  g0766(.A(new_n949_), .B1(new_n964_), .B2(new_n966_), .ZN(new_n967_));
  XNOR2_X1  g0767(.A(new_n708_), .B(KEYINPUT85), .ZN(new_n968_));
  OAI21_X1  g0768(.A(new_n945_), .B1(new_n967_), .B2(new_n968_), .ZN(new_n969_));
  NAND3_X1  g0769(.A1(new_n940_), .A2(new_n944_), .A3(new_n718_), .ZN(new_n970_));
  INV_X1    g0770(.A(KEYINPUT87), .ZN(new_n971_));
  AND2_X1   g0771(.A1(new_n240_), .A2(new_n778_), .ZN(new_n972_));
  OAI21_X1  g0772(.A(new_n777_), .B1(new_n210_), .B2(new_n509_), .ZN(new_n973_));
  OAI21_X1  g0773(.A(new_n720_), .B1(new_n972_), .B2(new_n973_), .ZN(new_n974_));
  INV_X1    g0774(.A(G311), .ZN(new_n975_));
  OAI22_X1  g0775(.A1(new_n732_), .A2(new_n975_), .B1(new_n734_), .B2(new_n593_), .ZN(new_n976_));
  AOI21_X1  g0776(.A(new_n976_), .B1(G283), .B2(new_n760_), .ZN(new_n977_));
  INV_X1    g0777(.A(G317), .ZN(new_n978_));
  OAI221_X1 g0778(.A(new_n977_), .B1(new_n214_), .B2(new_n754_), .C1(new_n978_), .C2(new_n847_), .ZN(new_n979_));
  AOI21_X1  g0779(.A(new_n299_), .B1(new_n759_), .B2(G294), .ZN(new_n980_));
  NAND2_X1  g0780(.A1(new_n832_), .A2(G97), .ZN(new_n981_));
  OAI211_X1 g0781(.A(new_n980_), .B(new_n981_), .C1(new_n611_), .C2(new_n745_), .ZN(new_n982_));
  NOR2_X1   g0782(.A1(new_n754_), .A2(new_n217_), .ZN(new_n983_));
  NOR2_X1   g0783(.A1(new_n740_), .A2(new_n838_), .ZN(new_n984_));
  INV_X1    g0784(.A(G143), .ZN(new_n985_));
  OAI22_X1  g0785(.A1(new_n732_), .A2(new_n985_), .B1(new_n734_), .B2(new_n837_), .ZN(new_n986_));
  NOR3_X1   g0786(.A1(new_n983_), .A2(new_n984_), .A3(new_n986_), .ZN(new_n987_));
  INV_X1    g0787(.A(G137), .ZN(new_n988_));
  OAI21_X1  g0788(.A(new_n987_), .B1(new_n988_), .B2(new_n847_), .ZN(new_n989_));
  AOI21_X1  g0789(.A(G33), .B1(new_n760_), .B2(G50), .ZN(new_n990_));
  OAI221_X1 g0790(.A(new_n990_), .B1(new_n265_), .B2(new_n745_), .C1(new_n202_), .C2(new_n747_), .ZN(new_n991_));
  OAI22_X1  g0791(.A1(new_n979_), .A2(new_n982_), .B1(new_n989_), .B2(new_n991_), .ZN(new_n992_));
  AOI21_X1  g0792(.A(new_n974_), .B1(new_n992_), .B2(new_n725_), .ZN(new_n993_));
  OAI21_X1  g0793(.A(new_n993_), .B1(new_n931_), .B2(new_n788_), .ZN(new_n994_));
  XOR2_X1   g0794(.A(new_n994_), .B(KEYINPUT86), .Z(new_n995_));
  AND3_X1   g0795(.A1(new_n970_), .A2(new_n971_), .A3(new_n995_), .ZN(new_n996_));
  AOI21_X1  g0796(.A(new_n971_), .B1(new_n970_), .B2(new_n995_), .ZN(new_n997_));
  OAI21_X1  g0797(.A(new_n969_), .B1(new_n996_), .B2(new_n997_), .ZN(new_n998_));
  XNOR2_X1  g0798(.A(new_n998_), .B(KEYINPUT88), .ZN(G387));
  NAND2_X1  g0799(.A1(new_n948_), .A2(new_n968_), .ZN(new_n1000_));
  XNOR2_X1  g0800(.A(new_n1000_), .B(KEYINPUT89), .ZN(new_n1001_));
  NAND3_X1  g0801(.A1(new_n1001_), .A2(new_n681_), .A3(new_n949_), .ZN(new_n1002_));
  NAND2_X1  g0802(.A1(new_n211_), .A2(new_n214_), .ZN(new_n1003_));
  NOR2_X1   g0803(.A1(new_n243_), .A2(new_n459_), .ZN(new_n1004_));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005_));
  NAND3_X1  g0805(.A1(new_n1005_), .A2(new_n328_), .A3(G58), .ZN(new_n1006_));
  OAI21_X1  g0806(.A(new_n778_), .B1(new_n684_), .B2(new_n1006_), .ZN(new_n1007_));
  OAI221_X1 g0807(.A(new_n1003_), .B1(new_n683_), .B2(new_n785_), .C1(new_n1004_), .C2(new_n1007_), .ZN(new_n1008_));
  AOI21_X1  g0808(.A(new_n721_), .B1(new_n1008_), .B2(new_n777_), .ZN(new_n1009_));
  OAI22_X1  g0809(.A1(new_n732_), .A2(new_n764_), .B1(new_n734_), .B2(new_n978_), .ZN(new_n1010_));
  XOR2_X1   g0810(.A(new_n1010_), .B(KEYINPUT91), .Z(new_n1011_));
  NOR2_X1   g0811(.A1(new_n741_), .A2(new_n593_), .ZN(new_n1012_));
  AOI211_X1 g0812(.A(new_n299_), .B(new_n1012_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n1013_));
  AOI22_X1  g0813(.A1(G116), .A2(new_n832_), .B1(new_n829_), .B2(G294), .ZN(new_n1014_));
  AOI22_X1  g0814(.A1(G283), .A2(new_n753_), .B1(new_n756_), .B2(G326), .ZN(new_n1015_));
  AND4_X1   g0815(.A1(new_n1011_), .A2(new_n1013_), .A3(new_n1014_), .A4(new_n1015_), .ZN(new_n1016_));
  AOI21_X1  g0816(.A(G33), .B1(new_n760_), .B2(G68), .ZN(new_n1017_));
  OAI211_X1 g0817(.A(new_n981_), .B(new_n1017_), .C1(new_n202_), .C2(new_n745_), .ZN(new_n1018_));
  AOI22_X1  g0818(.A1(G58), .A2(new_n759_), .B1(new_n733_), .B2(G159), .ZN(new_n1019_));
  OAI21_X1  g0819(.A(new_n1019_), .B1(new_n328_), .B2(new_n734_), .ZN(new_n1020_));
  AOI211_X1 g0820(.A(new_n1018_), .B(new_n1020_), .C1(G150), .C2(new_n756_), .ZN(new_n1021_));
  NAND2_X1  g0821(.A1(new_n753_), .A2(new_n394_), .ZN(new_n1022_));
  XNOR2_X1  g0822(.A(new_n1022_), .B(KEYINPUT90), .ZN(new_n1023_));
  AOI21_X1  g0823(.A(new_n1016_), .B1(new_n1021_), .B2(new_n1023_), .ZN(new_n1024_));
  NOR2_X1   g0824(.A1(new_n1024_), .A2(KEYINPUT92), .ZN(new_n1025_));
  NAND2_X1  g0825(.A1(new_n1024_), .A2(KEYINPUT92), .ZN(new_n1026_));
  NAND2_X1  g0826(.A1(new_n1026_), .A2(new_n725_), .ZN(new_n1027_));
  OAI221_X1 g0827(.A(new_n1009_), .B1(new_n1025_), .B2(new_n1027_), .C1(new_n668_), .C2(new_n788_), .ZN(new_n1028_));
  OAI21_X1  g0828(.A(new_n1028_), .B1(new_n948_), .B2(new_n716_), .ZN(new_n1029_));
  INV_X1    g0829(.A(new_n1029_), .ZN(new_n1030_));
  NAND2_X1  g0830(.A1(new_n1002_), .A2(new_n1030_), .ZN(G393));
  NAND2_X1  g0831(.A1(new_n964_), .A2(new_n966_), .ZN(new_n1032_));
  NAND2_X1  g0832(.A1(new_n1032_), .A2(new_n718_), .ZN(new_n1033_));
  OAI21_X1  g0833(.A(new_n777_), .B1(new_n224_), .B2(new_n210_), .ZN(new_n1034_));
  NOR2_X1   g0834(.A1(new_n247_), .A2(new_n779_), .ZN(new_n1035_));
  OAI21_X1  g0835(.A(new_n720_), .B1(new_n1034_), .B2(new_n1035_), .ZN(new_n1036_));
  NAND2_X1  g0836(.A1(new_n753_), .A2(G77), .ZN(new_n1037_));
  XOR2_X1   g0837(.A(new_n1037_), .B(KEYINPUT93), .Z(new_n1038_));
  INV_X1    g0838(.A(new_n1038_), .ZN(new_n1039_));
  OAI221_X1 g0839(.A(new_n299_), .B1(new_n732_), .B2(new_n837_), .C1(new_n219_), .C2(new_n747_), .ZN(new_n1040_));
  AOI21_X1  g0840(.A(new_n1040_), .B1(G68), .B2(new_n829_), .ZN(new_n1041_));
  NOR2_X1   g0841(.A1(new_n734_), .A2(new_n838_), .ZN(new_n1042_));
  OAI22_X1  g0842(.A1(new_n740_), .A2(new_n328_), .B1(new_n741_), .B2(new_n265_), .ZN(new_n1043_));
  AOI211_X1 g0843(.A(new_n1042_), .B(new_n1043_), .C1(G143), .C2(new_n756_), .ZN(new_n1044_));
  NAND3_X1  g0844(.A1(new_n1039_), .A2(new_n1041_), .A3(new_n1044_), .ZN(new_n1045_));
  OR2_X1    g0845(.A1(new_n1045_), .A2(KEYINPUT94), .ZN(new_n1046_));
  NOR2_X1   g0846(.A1(new_n732_), .A2(new_n978_), .ZN(new_n1047_));
  OAI22_X1  g0847(.A1(new_n740_), .A2(new_n593_), .B1(new_n734_), .B2(new_n975_), .ZN(new_n1048_));
  AOI211_X1 g0848(.A(new_n1047_), .B(new_n1048_), .C1(G322), .C2(new_n756_), .ZN(new_n1049_));
  AOI211_X1 g0849(.A(new_n299_), .B(new_n748_), .C1(G294), .C2(new_n760_), .ZN(new_n1050_));
  NAND2_X1  g0850(.A1(new_n829_), .A2(G283), .ZN(new_n1051_));
  NAND2_X1  g0851(.A1(new_n753_), .A2(G116), .ZN(new_n1052_));
  NAND4_X1  g0852(.A1(new_n1049_), .A2(new_n1050_), .A3(new_n1051_), .A4(new_n1052_), .ZN(new_n1053_));
  NAND2_X1  g0853(.A1(new_n1045_), .A2(KEYINPUT94), .ZN(new_n1054_));
  NAND3_X1  g0854(.A1(new_n1046_), .A2(new_n1053_), .A3(new_n1054_), .ZN(new_n1055_));
  AOI21_X1  g0855(.A(new_n1036_), .B1(new_n1055_), .B2(new_n725_), .ZN(new_n1056_));
  OAI21_X1  g0856(.A(new_n1056_), .B1(new_n922_), .B2(new_n788_), .ZN(new_n1057_));
  NAND3_X1  g0857(.A1(new_n965_), .A2(new_n949_), .A3(new_n961_), .ZN(new_n1058_));
  NAND2_X1  g0858(.A1(new_n1058_), .A2(new_n681_), .ZN(new_n1059_));
  OAI211_X1 g0859(.A(new_n1033_), .B(new_n1057_), .C1(new_n967_), .C2(new_n1059_), .ZN(G390));
  NAND3_X1  g0860(.A1(new_n445_), .A2(new_n672_), .A3(new_n698_), .ZN(new_n1061_));
  NAND3_X1  g0861(.A1(new_n905_), .A2(new_n1061_), .A3(new_n650_), .ZN(new_n1062_));
  XNOR2_X1  g0862(.A(new_n1062_), .B(KEYINPUT100), .ZN(new_n1063_));
  INV_X1    g0863(.A(KEYINPUT99), .ZN(new_n1064_));
  NAND4_X1  g0864(.A1(new_n696_), .A2(G330), .A3(new_n697_), .A4(new_n801_), .ZN(new_n1065_));
  NAND2_X1  g0865(.A1(new_n1065_), .A2(KEYINPUT97), .ZN(new_n1066_));
  AND3_X1   g0866(.A1(new_n890_), .A2(new_n883_), .A3(new_n892_), .ZN(new_n1067_));
  AOI21_X1  g0867(.A(new_n883_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n1068_));
  OAI21_X1  g0868(.A(new_n1066_), .B1(new_n1067_), .B2(new_n1068_), .ZN(new_n1069_));
  NOR2_X1   g0869(.A1(new_n1065_), .A2(KEYINPUT97), .ZN(new_n1070_));
  OAI21_X1  g0870(.A(KEYINPUT98), .B1(new_n1069_), .B2(new_n1070_), .ZN(new_n1071_));
  AOI21_X1  g0871(.A(new_n881_), .B1(new_n389_), .B2(new_n877_), .ZN(new_n1072_));
  NAND2_X1  g0872(.A1(new_n893_), .A2(new_n1072_), .ZN(new_n1073_));
  NAND3_X1  g0873(.A1(new_n890_), .A2(new_n883_), .A3(new_n892_), .ZN(new_n1074_));
  NAND2_X1  g0874(.A1(new_n1073_), .A2(new_n1074_), .ZN(new_n1075_));
  OR2_X1    g0875(.A1(new_n1065_), .A2(KEYINPUT97), .ZN(new_n1076_));
  INV_X1    g0876(.A(KEYINPUT98), .ZN(new_n1077_));
  NAND4_X1  g0877(.A1(new_n1075_), .A2(new_n1076_), .A3(new_n1077_), .A4(new_n1066_), .ZN(new_n1078_));
  NAND2_X1  g0878(.A1(new_n1071_), .A2(new_n1078_), .ZN(new_n1079_));
  NAND4_X1  g0879(.A1(new_n805_), .A2(new_n672_), .A3(new_n696_), .A4(new_n697_), .ZN(new_n1080_));
  NAND2_X1  g0880(.A1(new_n1072_), .A2(KEYINPUT96), .ZN(new_n1081_));
  AND3_X1   g0881(.A1(new_n890_), .A2(new_n892_), .A3(new_n1081_), .ZN(new_n1082_));
  AOI21_X1  g0882(.A(new_n1081_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n1083_));
  NOR3_X1   g0883(.A1(new_n1080_), .A2(new_n1082_), .A3(new_n1083_), .ZN(new_n1084_));
  INV_X1    g0884(.A(new_n1084_), .ZN(new_n1085_));
  AOI21_X1  g0885(.A(new_n1064_), .B1(new_n1079_), .B2(new_n1085_), .ZN(new_n1086_));
  AOI211_X1 g0886(.A(KEYINPUT99), .B(new_n1084_), .C1(new_n1071_), .C2(new_n1078_), .ZN(new_n1087_));
  OAI21_X1  g0887(.A(new_n1063_), .B1(new_n1086_), .B2(new_n1087_), .ZN(new_n1088_));
  OR2_X1    g0888(.A1(new_n1065_), .A2(new_n1072_), .ZN(new_n1089_));
  NAND4_X1  g0889(.A1(new_n644_), .A2(new_n659_), .A3(new_n801_), .A4(new_n883_), .ZN(new_n1090_));
  OAI21_X1  g0890(.A(KEYINPUT95), .B1(new_n1072_), .B2(new_n892_), .ZN(new_n1091_));
  INV_X1    g0891(.A(KEYINPUT95), .ZN(new_n1092_));
  NAND3_X1  g0892(.A1(new_n883_), .A2(new_n1092_), .A3(new_n891_), .ZN(new_n1093_));
  AOI21_X1  g0893(.A(new_n900_), .B1(new_n1091_), .B2(new_n1093_), .ZN(new_n1094_));
  AND3_X1   g0894(.A1(new_n1090_), .A2(new_n1094_), .A3(new_n876_), .ZN(new_n1095_));
  AOI21_X1  g0895(.A(new_n876_), .B1(new_n1090_), .B2(new_n1094_), .ZN(new_n1096_));
  OAI21_X1  g0896(.A(new_n1089_), .B1(new_n1095_), .B2(new_n1096_), .ZN(new_n1097_));
  INV_X1    g0897(.A(new_n876_), .ZN(new_n1098_));
  INV_X1    g0898(.A(new_n900_), .ZN(new_n1099_));
  NOR3_X1   g0899(.A1(new_n1072_), .A2(new_n892_), .A3(KEYINPUT95), .ZN(new_n1100_));
  AOI21_X1  g0900(.A(new_n1092_), .B1(new_n883_), .B2(new_n891_), .ZN(new_n1101_));
  OAI21_X1  g0901(.A(new_n1099_), .B1(new_n1100_), .B2(new_n1101_), .ZN(new_n1102_));
  NOR2_X1   g0902(.A1(new_n890_), .A2(new_n1072_), .ZN(new_n1103_));
  OAI21_X1  g0903(.A(new_n1098_), .B1(new_n1102_), .B2(new_n1103_), .ZN(new_n1104_));
  NAND3_X1  g0904(.A1(new_n1090_), .A2(new_n1094_), .A3(new_n876_), .ZN(new_n1105_));
  NOR2_X1   g0905(.A1(new_n1065_), .A2(new_n1072_), .ZN(new_n1106_));
  NAND3_X1  g0906(.A1(new_n1104_), .A2(new_n1105_), .A3(new_n1106_), .ZN(new_n1107_));
  NAND2_X1  g0907(.A1(new_n1097_), .A2(new_n1107_), .ZN(new_n1108_));
  INV_X1    g0908(.A(new_n1108_), .ZN(new_n1109_));
  NAND2_X1  g0909(.A1(new_n1088_), .A2(new_n1109_), .ZN(new_n1110_));
  OAI211_X1 g0910(.A(new_n1108_), .B(new_n1063_), .C1(new_n1086_), .C2(new_n1087_), .ZN(new_n1111_));
  NAND3_X1  g0911(.A1(new_n1110_), .A2(new_n681_), .A3(new_n1111_), .ZN(new_n1112_));
  NOR3_X1   g0912(.A1(new_n1095_), .A2(new_n1089_), .A3(new_n1096_), .ZN(new_n1113_));
  AOI21_X1  g0913(.A(new_n1106_), .B1(new_n1104_), .B2(new_n1105_), .ZN(new_n1114_));
  OAI21_X1  g0914(.A(new_n718_), .B1(new_n1113_), .B2(new_n1114_), .ZN(new_n1115_));
  INV_X1    g0915(.A(KEYINPUT105), .ZN(new_n1116_));
  NAND2_X1  g0916(.A1(new_n1098_), .A2(new_n773_), .ZN(new_n1117_));
  XOR2_X1   g0917(.A(new_n1117_), .B(KEYINPUT104), .Z(new_n1118_));
  OAI22_X1  g0918(.A1(new_n732_), .A2(new_n769_), .B1(new_n741_), .B2(new_n224_), .ZN(new_n1119_));
  OAI22_X1  g0919(.A1(new_n740_), .A2(new_n577_), .B1(new_n734_), .B2(new_n611_), .ZN(new_n1120_));
  NOR4_X1   g0920(.A1(new_n1038_), .A2(new_n746_), .A3(new_n1119_), .A4(new_n1120_), .ZN(new_n1121_));
  XNOR2_X1  g0921(.A(new_n1121_), .B(KEYINPUT102), .ZN(new_n1122_));
  NAND2_X1  g0922(.A1(new_n756_), .A2(G294), .ZN(new_n1123_));
  XOR2_X1   g0923(.A(new_n1123_), .B(KEYINPUT103), .Z(new_n1124_));
  OAI21_X1  g0924(.A(G33), .B1(new_n747_), .B2(new_n217_), .ZN(new_n1125_));
  NOR3_X1   g0925(.A1(new_n1122_), .A2(new_n1124_), .A3(new_n1125_), .ZN(new_n1126_));
  AOI22_X1  g0926(.A1(G128), .A2(new_n733_), .B1(new_n759_), .B2(G137), .ZN(new_n1127_));
  OAI221_X1 g0927(.A(new_n1127_), .B1(new_n985_), .B2(new_n741_), .C1(new_n838_), .C2(new_n754_), .ZN(new_n1128_));
  NAND2_X1  g0928(.A1(new_n756_), .A2(G125), .ZN(new_n1129_));
  XNOR2_X1  g0929(.A(new_n1129_), .B(KEYINPUT101), .ZN(new_n1130_));
  AOI21_X1  g0930(.A(G33), .B1(new_n735_), .B2(G132), .ZN(new_n1131_));
  OAI221_X1 g0931(.A(new_n1131_), .B1(new_n745_), .B2(new_n837_), .C1(new_n328_), .C2(new_n747_), .ZN(new_n1132_));
  NOR3_X1   g0932(.A1(new_n1128_), .A2(new_n1130_), .A3(new_n1132_), .ZN(new_n1133_));
  OAI21_X1  g0933(.A(new_n725_), .B1(new_n1126_), .B2(new_n1133_), .ZN(new_n1134_));
  OAI211_X1 g0934(.A(new_n1134_), .B(new_n720_), .C1(G58), .C2(new_n825_), .ZN(new_n1135_));
  NOR2_X1   g0935(.A1(new_n1118_), .A2(new_n1135_), .ZN(new_n1136_));
  INV_X1    g0936(.A(new_n1136_), .ZN(new_n1137_));
  NAND3_X1  g0937(.A1(new_n1115_), .A2(new_n1116_), .A3(new_n1137_), .ZN(new_n1138_));
  AOI21_X1  g0938(.A(new_n717_), .B1(new_n1097_), .B2(new_n1107_), .ZN(new_n1139_));
  OAI21_X1  g0939(.A(KEYINPUT105), .B1(new_n1139_), .B2(new_n1136_), .ZN(new_n1140_));
  NAND2_X1  g0940(.A1(new_n1138_), .A2(new_n1140_), .ZN(new_n1141_));
  NAND2_X1  g0941(.A1(new_n1112_), .A2(new_n1141_), .ZN(G378));
  NOR2_X1   g0942(.A1(new_n901_), .A2(KEYINPUT106), .ZN(new_n1143_));
  INV_X1    g0943(.A(KEYINPUT106), .ZN(new_n1144_));
  AOI21_X1  g0944(.A(new_n1144_), .B1(new_n876_), .B2(new_n900_), .ZN(new_n1145_));
  NOR2_X1   g0945(.A1(new_n1143_), .A2(new_n1145_), .ZN(new_n1146_));
  NAND2_X1  g0946(.A1(new_n331_), .A2(new_n860_), .ZN(new_n1147_));
  XNOR2_X1  g0947(.A(new_n346_), .B(new_n1147_), .ZN(new_n1148_));
  NOR2_X1   g0948(.A1(new_n1146_), .A2(new_n1148_), .ZN(new_n1149_));
  NOR2_X1   g0949(.A1(new_n902_), .A2(new_n897_), .ZN(new_n1150_));
  NAND2_X1  g0950(.A1(new_n1149_), .A2(new_n1150_), .ZN(new_n1151_));
  INV_X1    g0951(.A(new_n904_), .ZN(new_n1152_));
  INV_X1    g0952(.A(new_n1148_), .ZN(new_n1153_));
  OAI21_X1  g0953(.A(new_n1151_), .B1(new_n1152_), .B2(new_n1153_), .ZN(new_n1154_));
  NAND3_X1  g0954(.A1(new_n698_), .A2(new_n885_), .A3(new_n672_), .ZN(new_n1155_));
  NAND2_X1  g0955(.A1(new_n1154_), .A2(new_n1155_), .ZN(new_n1156_));
  INV_X1    g0956(.A(KEYINPUT107), .ZN(new_n1157_));
  AOI22_X1  g0957(.A1(new_n904_), .A2(new_n1148_), .B1(new_n1150_), .B2(new_n1149_), .ZN(new_n1158_));
  INV_X1    g0958(.A(new_n1155_), .ZN(new_n1159_));
  AOI21_X1  g0959(.A(new_n1157_), .B1(new_n1158_), .B2(new_n1159_), .ZN(new_n1160_));
  NAND2_X1  g0960(.A1(new_n1156_), .A2(new_n1160_), .ZN(new_n1161_));
  NAND3_X1  g0961(.A1(new_n1154_), .A2(new_n1157_), .A3(new_n1155_), .ZN(new_n1162_));
  NAND3_X1  g0962(.A1(new_n1161_), .A2(new_n681_), .A3(new_n1162_), .ZN(new_n1163_));
  INV_X1    g0963(.A(new_n1163_), .ZN(new_n1164_));
  NAND2_X1  g0964(.A1(new_n1111_), .A2(new_n1063_), .ZN(new_n1165_));
  NAND3_X1  g0965(.A1(new_n1164_), .A2(KEYINPUT108), .A3(new_n1165_), .ZN(new_n1166_));
  INV_X1    g0966(.A(KEYINPUT108), .ZN(new_n1167_));
  INV_X1    g0967(.A(new_n1063_), .ZN(new_n1168_));
  NAND2_X1  g0968(.A1(new_n1079_), .A2(new_n1085_), .ZN(new_n1169_));
  NAND2_X1  g0969(.A1(new_n1169_), .A2(KEYINPUT99), .ZN(new_n1170_));
  NAND3_X1  g0970(.A1(new_n1079_), .A2(new_n1064_), .A3(new_n1085_), .ZN(new_n1171_));
  NAND2_X1  g0971(.A1(new_n1170_), .A2(new_n1171_), .ZN(new_n1172_));
  AOI21_X1  g0972(.A(new_n1168_), .B1(new_n1172_), .B2(new_n1108_), .ZN(new_n1173_));
  OAI21_X1  g0973(.A(new_n1167_), .B1(new_n1173_), .B2(new_n1163_), .ZN(new_n1174_));
  AOI22_X1  g0974(.A1(new_n733_), .A2(G116), .B1(new_n735_), .B2(G107), .ZN(new_n1175_));
  OAI221_X1 g0975(.A(new_n1175_), .B1(new_n224_), .B2(new_n740_), .C1(new_n509_), .C2(new_n741_), .ZN(new_n1176_));
  XNOR2_X1  g0976(.A(new_n1176_), .B(KEYINPUT111), .ZN(new_n1177_));
  NAND2_X1  g0977(.A1(new_n455_), .A2(G33), .ZN(new_n1178_));
  XNOR2_X1  g0978(.A(new_n1178_), .B(KEYINPUT112), .ZN(new_n1179_));
  AOI21_X1  g0979(.A(new_n1179_), .B1(new_n829_), .B2(G77), .ZN(new_n1180_));
  OAI21_X1  g0980(.A(new_n1180_), .B1(new_n265_), .B2(new_n747_), .ZN(new_n1181_));
  AOI211_X1 g0981(.A(new_n983_), .B(new_n1181_), .C1(G283), .C2(new_n756_), .ZN(new_n1182_));
  NAND2_X1  g0982(.A1(new_n1177_), .A2(new_n1182_), .ZN(new_n1183_));
  OAI211_X1 g0983(.A(new_n1179_), .B(new_n328_), .C1(G33), .C2(G41), .ZN(new_n1184_));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n760_), .C2(G137), .ZN(new_n1185_));
  OAI221_X1 g0985(.A(new_n1185_), .B1(new_n985_), .B2(new_n745_), .C1(new_n838_), .C2(new_n747_), .ZN(new_n1186_));
  INV_X1    g0986(.A(G128), .ZN(new_n1187_));
  OAI22_X1  g0987(.A1(new_n740_), .A2(new_n848_), .B1(new_n734_), .B2(new_n1187_), .ZN(new_n1188_));
  AOI21_X1  g0988(.A(new_n1188_), .B1(G125), .B2(new_n733_), .ZN(new_n1189_));
  NAND2_X1  g0989(.A1(new_n756_), .A2(G124), .ZN(new_n1190_));
  OAI211_X1 g0990(.A(new_n1189_), .B(new_n1190_), .C1(new_n837_), .C2(new_n754_), .ZN(new_n1191_));
  OAI211_X1 g0991(.A(new_n1183_), .B(new_n1184_), .C1(new_n1186_), .C2(new_n1191_), .ZN(new_n1192_));
  INV_X1    g0992(.A(KEYINPUT113), .ZN(new_n1193_));
  OR2_X1    g0993(.A1(new_n1192_), .A2(new_n1193_), .ZN(new_n1194_));
  NAND2_X1  g0994(.A1(new_n1192_), .A2(new_n1193_), .ZN(new_n1195_));
  NAND3_X1  g0995(.A1(new_n1194_), .A2(new_n725_), .A3(new_n1195_), .ZN(new_n1196_));
  AOI21_X1  g0996(.A(new_n721_), .B1(new_n328_), .B2(new_n824_), .ZN(new_n1197_));
  OAI211_X1 g0997(.A(new_n1196_), .B(new_n1197_), .C1(new_n1153_), .C2(new_n775_), .ZN(new_n1198_));
  AOI221_X4 g0998(.A(new_n1155_), .B1(new_n1149_), .B2(new_n1150_), .C1(new_n904_), .C2(new_n1148_), .ZN(new_n1199_));
  AOI21_X1  g0999(.A(new_n896_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n1200_));
  NOR3_X1   g1000(.A1(new_n902_), .A2(KEYINPUT74), .A3(new_n897_), .ZN(new_n1201_));
  NOR2_X1   g1001(.A1(new_n1200_), .A2(new_n1201_), .ZN(new_n1202_));
  INV_X1    g1002(.A(KEYINPUT110), .ZN(new_n1203_));
  NAND4_X1  g1003(.A1(new_n1202_), .A2(new_n1203_), .A3(new_n901_), .A4(new_n1153_), .ZN(new_n1204_));
  OAI21_X1  g1004(.A(KEYINPUT110), .B1(new_n904_), .B2(new_n1148_), .ZN(new_n1205_));
  OAI211_X1 g1005(.A(new_n899_), .B(new_n903_), .C1(new_n1145_), .C2(new_n1143_), .ZN(new_n1206_));
  NAND2_X1  g1006(.A1(new_n1206_), .A2(new_n1148_), .ZN(new_n1207_));
  NAND3_X1  g1007(.A1(new_n1204_), .A2(new_n1205_), .A3(new_n1207_), .ZN(new_n1208_));
  XOR2_X1   g1008(.A(new_n1155_), .B(KEYINPUT109), .Z(new_n1209_));
  AOI21_X1  g1009(.A(new_n1199_), .B1(new_n1208_), .B2(new_n1209_), .ZN(new_n1210_));
  OAI21_X1  g1010(.A(new_n1198_), .B1(new_n1210_), .B2(new_n717_), .ZN(new_n1211_));
  INV_X1    g1011(.A(new_n1211_), .ZN(new_n1212_));
  NAND3_X1  g1012(.A1(new_n1166_), .A2(new_n1174_), .A3(new_n1212_), .ZN(G375));
  NAND3_X1  g1013(.A1(new_n1168_), .A2(new_n1170_), .A3(new_n1171_), .ZN(new_n1214_));
  NAND3_X1  g1014(.A1(new_n1214_), .A2(new_n1088_), .A3(new_n681_), .ZN(new_n1215_));
  XOR2_X1   g1015(.A(new_n1215_), .B(KEYINPUT114), .Z(new_n1216_));
  OAI221_X1 g1016(.A(G33), .B1(new_n740_), .B2(new_n611_), .C1(new_n202_), .C2(new_n747_), .ZN(new_n1217_));
  AOI22_X1  g1017(.A1(new_n733_), .A2(G294), .B1(new_n760_), .B2(new_n576_), .ZN(new_n1218_));
  OAI221_X1 g1018(.A(new_n1218_), .B1(new_n769_), .B2(new_n734_), .C1(new_n593_), .C2(new_n847_), .ZN(new_n1219_));
  AOI211_X1 g1019(.A(new_n1217_), .B(new_n1219_), .C1(G97), .C2(new_n829_), .ZN(new_n1220_));
  NAND2_X1  g1020(.A1(new_n829_), .A2(G159), .ZN(new_n1221_));
  XNOR2_X1  g1021(.A(new_n1221_), .B(KEYINPUT115), .ZN(new_n1222_));
  AOI22_X1  g1022(.A1(new_n733_), .A2(G132), .B1(new_n760_), .B2(G150), .ZN(new_n1223_));
  OAI21_X1  g1023(.A(new_n1223_), .B1(new_n988_), .B2(new_n734_), .ZN(new_n1224_));
  OAI221_X1 g1024(.A(new_n299_), .B1(new_n740_), .B2(new_n985_), .C1(new_n265_), .C2(new_n747_), .ZN(new_n1225_));
  OAI22_X1  g1025(.A1(new_n328_), .A2(new_n754_), .B1(new_n847_), .B2(new_n1187_), .ZN(new_n1226_));
  NOR3_X1   g1026(.A1(new_n1224_), .A2(new_n1225_), .A3(new_n1226_), .ZN(new_n1227_));
  AOI22_X1  g1027(.A1(new_n1220_), .A2(new_n1023_), .B1(new_n1222_), .B2(new_n1227_), .ZN(new_n1228_));
  OAI221_X1 g1028(.A(new_n720_), .B1(G68), .B2(new_n825_), .C1(new_n1228_), .C2(new_n726_), .ZN(new_n1229_));
  AOI21_X1  g1029(.A(new_n1229_), .B1(new_n773_), .B2(new_n1072_), .ZN(new_n1230_));
  AOI21_X1  g1030(.A(new_n1230_), .B1(new_n1172_), .B2(new_n718_), .ZN(new_n1231_));
  NAND2_X1  g1031(.A1(new_n1216_), .A2(new_n1231_), .ZN(G381));
  INV_X1    g1032(.A(G396), .ZN(new_n1233_));
  NAND3_X1  g1033(.A1(new_n1002_), .A2(new_n1233_), .A3(new_n1030_), .ZN(new_n1234_));
  OR3_X1    g1034(.A1(G390), .A2(G384), .A3(new_n1234_), .ZN(new_n1235_));
  OR3_X1    g1035(.A1(new_n1235_), .A2(G378), .A3(G381), .ZN(new_n1236_));
  OR3_X1    g1036(.A1(new_n1236_), .A2(G387), .A3(G375), .ZN(G407));
  OR3_X1    g1037(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1238_));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238_), .ZN(G409));
  NAND2_X1  g1039(.A1(new_n1215_), .A2(new_n1231_), .ZN(new_n1240_));
  INV_X1    g1040(.A(G384), .ZN(new_n1241_));
  NAND2_X1  g1041(.A1(new_n1240_), .A2(new_n1241_), .ZN(new_n1242_));
  NAND3_X1  g1042(.A1(new_n1215_), .A2(G384), .A3(new_n1231_), .ZN(new_n1243_));
  NAND2_X1  g1043(.A1(new_n1242_), .A2(new_n1243_), .ZN(new_n1244_));
  NAND3_X1  g1044(.A1(new_n657_), .A2(G213), .A3(G2897), .ZN(new_n1245_));
  NOR2_X1   g1045(.A1(new_n1244_), .A2(new_n1245_), .ZN(new_n1246_));
  OR2_X1    g1046(.A1(new_n1246_), .A2(KEYINPUT125), .ZN(new_n1247_));
  NAND2_X1  g1047(.A1(new_n1246_), .A2(KEYINPUT125), .ZN(new_n1248_));
  NAND2_X1  g1048(.A1(new_n657_), .A2(G213), .ZN(new_n1249_));
  INV_X1    g1049(.A(KEYINPUT116), .ZN(new_n1250_));
  AND3_X1   g1050(.A1(new_n1138_), .A2(new_n1140_), .A3(new_n1250_), .ZN(new_n1251_));
  AOI21_X1  g1051(.A(new_n1250_), .B1(new_n1138_), .B2(new_n1140_), .ZN(new_n1252_));
  NOR2_X1   g1052(.A1(new_n1251_), .A2(new_n1252_), .ZN(new_n1253_));
  NAND3_X1  g1053(.A1(new_n1112_), .A2(KEYINPUT117), .A3(new_n1253_), .ZN(new_n1254_));
  INV_X1    g1054(.A(new_n1254_), .ZN(new_n1255_));
  NAND3_X1  g1055(.A1(new_n1161_), .A2(new_n1168_), .A3(new_n1162_), .ZN(new_n1256_));
  OAI21_X1  g1056(.A(new_n1256_), .B1(new_n1111_), .B2(new_n1210_), .ZN(new_n1257_));
  AOI21_X1  g1057(.A(new_n1211_), .B1(new_n1257_), .B2(new_n681_), .ZN(new_n1258_));
  AOI21_X1  g1058(.A(KEYINPUT117), .B1(new_n1112_), .B2(new_n1253_), .ZN(new_n1259_));
  NOR3_X1   g1059(.A1(new_n1255_), .A2(new_n1258_), .A3(new_n1259_), .ZN(new_n1260_));
  NAND4_X1  g1060(.A1(G378), .A2(new_n1166_), .A3(new_n1212_), .A4(new_n1174_), .ZN(new_n1261_));
  INV_X1    g1061(.A(new_n1261_), .ZN(new_n1262_));
  OAI21_X1  g1062(.A(new_n1249_), .B1(new_n1260_), .B2(new_n1262_), .ZN(new_n1263_));
  INV_X1    g1063(.A(KEYINPUT119), .ZN(new_n1264_));
  INV_X1    g1064(.A(new_n1245_), .ZN(new_n1265_));
  OAI21_X1  g1065(.A(new_n1264_), .B1(new_n1244_), .B2(new_n1265_), .ZN(new_n1266_));
  NAND4_X1  g1066(.A1(new_n1242_), .A2(KEYINPUT119), .A3(new_n1243_), .A4(new_n1245_), .ZN(new_n1267_));
  NAND2_X1  g1067(.A1(new_n1266_), .A2(new_n1267_), .ZN(new_n1268_));
  OAI211_X1 g1068(.A(new_n1247_), .B(new_n1248_), .C1(new_n1263_), .C2(new_n1268_), .ZN(new_n1269_));
  OR2_X1    g1069(.A1(new_n1269_), .A2(KEYINPUT126), .ZN(new_n1270_));
  NAND2_X1  g1070(.A1(new_n1244_), .A2(new_n1245_), .ZN(new_n1271_));
  AND3_X1   g1071(.A1(new_n1161_), .A2(new_n1168_), .A3(new_n1162_), .ZN(new_n1272_));
  NOR2_X1   g1072(.A1(new_n1111_), .A2(new_n1210_), .ZN(new_n1273_));
  OAI21_X1  g1073(.A(new_n681_), .B1(new_n1272_), .B2(new_n1273_), .ZN(new_n1274_));
  NAND2_X1  g1074(.A1(new_n1274_), .A2(new_n1212_), .ZN(new_n1275_));
  AOI21_X1  g1075(.A(new_n1108_), .B1(new_n1172_), .B2(new_n1063_), .ZN(new_n1276_));
  NAND2_X1  g1076(.A1(new_n1111_), .A2(new_n681_), .ZN(new_n1277_));
  OAI21_X1  g1077(.A(new_n1253_), .B1(new_n1276_), .B2(new_n1277_), .ZN(new_n1278_));
  INV_X1    g1078(.A(KEYINPUT117), .ZN(new_n1279_));
  NAND2_X1  g1079(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1280_));
  NAND3_X1  g1080(.A1(new_n1275_), .A2(new_n1254_), .A3(new_n1280_), .ZN(new_n1281_));
  NAND2_X1  g1081(.A1(new_n1281_), .A2(new_n1261_), .ZN(new_n1282_));
  AOI21_X1  g1082(.A(new_n1271_), .B1(new_n1282_), .B2(new_n1249_), .ZN(new_n1283_));
  AOI22_X1  g1083(.A1(new_n1281_), .A2(new_n1261_), .B1(G213), .B2(new_n657_), .ZN(new_n1284_));
  INV_X1    g1084(.A(new_n1243_), .ZN(new_n1285_));
  AOI21_X1  g1085(.A(G384), .B1(new_n1231_), .B2(new_n1215_), .ZN(new_n1286_));
  OAI21_X1  g1086(.A(new_n1265_), .B1(new_n1285_), .B2(new_n1286_), .ZN(new_n1287_));
  INV_X1    g1087(.A(KEYINPUT118), .ZN(new_n1288_));
  NAND2_X1  g1088(.A1(new_n1287_), .A2(new_n1288_), .ZN(new_n1289_));
  NAND3_X1  g1089(.A1(new_n1244_), .A2(KEYINPUT118), .A3(new_n1265_), .ZN(new_n1290_));
  AND2_X1   g1090(.A1(new_n1289_), .A2(new_n1290_), .ZN(new_n1291_));
  AOI21_X1  g1091(.A(new_n1283_), .B1(new_n1284_), .B2(new_n1291_), .ZN(new_n1292_));
  NAND2_X1  g1092(.A1(new_n1269_), .A2(KEYINPUT126), .ZN(new_n1293_));
  INV_X1    g1093(.A(G390), .ZN(new_n1294_));
  NAND2_X1  g1094(.A1(new_n998_), .A2(new_n1294_), .ZN(new_n1295_));
  OAI211_X1 g1095(.A(G390), .B(new_n969_), .C1(new_n997_), .C2(new_n996_), .ZN(new_n1296_));
  NAND2_X1  g1096(.A1(new_n1295_), .A2(new_n1296_), .ZN(new_n1297_));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298_));
  NAND2_X1  g1098(.A1(new_n1298_), .A2(new_n1234_), .ZN(new_n1299_));
  INV_X1    g1099(.A(new_n1299_), .ZN(new_n1300_));
  XNOR2_X1  g1100(.A(new_n1297_), .B(new_n1300_), .ZN(new_n1301_));
  NAND4_X1  g1101(.A1(new_n1270_), .A2(new_n1292_), .A3(new_n1293_), .A4(new_n1301_), .ZN(new_n1302_));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303_));
  NAND3_X1  g1103(.A1(new_n1242_), .A2(new_n1243_), .A3(new_n1265_), .ZN(new_n1304_));
  XOR2_X1   g1104(.A(new_n1304_), .B(KEYINPUT121), .Z(new_n1305_));
  OAI21_X1  g1105(.A(KEYINPUT120), .B1(new_n1263_), .B2(new_n1268_), .ZN(new_n1306_));
  INV_X1    g1106(.A(KEYINPUT120), .ZN(new_n1307_));
  NAND4_X1  g1107(.A1(new_n1284_), .A2(new_n1307_), .A3(new_n1266_), .A4(new_n1267_), .ZN(new_n1308_));
  NAND4_X1  g1108(.A1(new_n1292_), .A2(new_n1305_), .A3(new_n1306_), .A4(new_n1308_), .ZN(new_n1309_));
  NAND3_X1  g1109(.A1(new_n1298_), .A2(KEYINPUT123), .A3(new_n1234_), .ZN(new_n1310_));
  AOI22_X1  g1110(.A1(new_n1295_), .A2(new_n1296_), .B1(new_n1310_), .B2(KEYINPUT122), .ZN(new_n1311_));
  NAND3_X1  g1111(.A1(new_n1295_), .A2(new_n1296_), .A3(KEYINPUT122), .ZN(new_n1312_));
  NAND2_X1  g1112(.A1(new_n1312_), .A2(KEYINPUT123), .ZN(new_n1313_));
  AOI21_X1  g1113(.A(new_n1311_), .B1(new_n1313_), .B2(new_n1299_), .ZN(new_n1314_));
  AOI21_X1  g1114(.A(new_n1303_), .B1(new_n1309_), .B2(new_n1314_), .ZN(new_n1315_));
  NAND2_X1  g1115(.A1(new_n1306_), .A2(new_n1308_), .ZN(new_n1316_));
  NAND4_X1  g1116(.A1(new_n1282_), .A2(new_n1289_), .A3(new_n1249_), .A4(new_n1290_), .ZN(new_n1317_));
  OAI211_X1 g1117(.A(new_n1305_), .B(new_n1317_), .C1(new_n1284_), .C2(new_n1271_), .ZN(new_n1318_));
  OAI211_X1 g1118(.A(new_n1303_), .B(new_n1314_), .C1(new_n1316_), .C2(new_n1318_), .ZN(new_n1319_));
  INV_X1    g1119(.A(new_n1319_), .ZN(new_n1320_));
  OAI21_X1  g1120(.A(new_n1302_), .B1(new_n1315_), .B2(new_n1320_), .ZN(G405));
  NAND2_X1  g1121(.A1(new_n1261_), .A2(KEYINPUT127), .ZN(new_n1322_));
  NAND2_X1  g1122(.A1(new_n1322_), .A2(new_n1244_), .ZN(new_n1323_));
  NAND2_X1  g1123(.A1(new_n1314_), .A2(new_n1323_), .ZN(new_n1324_));
  AOI21_X1  g1124(.A(new_n1300_), .B1(new_n1312_), .B2(KEYINPUT123), .ZN(new_n1325_));
  OAI211_X1 g1125(.A(new_n1244_), .B(new_n1322_), .C1(new_n1325_), .C2(new_n1311_), .ZN(new_n1326_));
  NAND2_X1  g1126(.A1(new_n1324_), .A2(new_n1326_), .ZN(new_n1327_));
  XNOR2_X1  g1127(.A(G375), .B(G378), .ZN(new_n1328_));
  INV_X1    g1128(.A(new_n1328_), .ZN(new_n1329_));
  NAND2_X1  g1129(.A1(new_n1327_), .A2(new_n1329_), .ZN(new_n1330_));
  NAND3_X1  g1130(.A1(new_n1324_), .A2(new_n1328_), .A3(new_n1326_), .ZN(new_n1331_));
  NAND2_X1  g1131(.A1(new_n1330_), .A2(new_n1331_), .ZN(G402));
endmodule


