//Secret key is'0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_c5315" written by ABC on Sun Nov 20 19:50:27 2022

module locked_c5315 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G1, G4, G11, G14, G17, G20, G23, G24, G25,
    G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64,
    G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94,
    G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161,
    G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197,
    G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241,
    G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281,
    G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324,
    G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372,
    G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479,
    G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562,
    G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546,
    G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091,
    G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G1, G4, G11, G14, G17, G20, G23,
    G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54,
    G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88,
    G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116,
    G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130,
    G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155,
    G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191,
    G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233,
    G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273,
    G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316,
    G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366,
    G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457,
    G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559,
    G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173,
    G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090,
    G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_n444_, new_n449_, new_n451_, new_n461_, new_n469_, new_n470_,
    new_n472_, new_n476_, new_n477_, new_n478_, new_n480_, new_n481_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n490_, new_n491_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1114_, new_n1115_, new_n1116_, new_n1118_,
    new_n1119_, new_n1120_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1128_, new_n1129_, new_n1130_, new_n1132_, new_n1133_,
    new_n1134_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1213_, new_n1214_, new_n1215_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1227_,
    new_n1228_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1235_,
    new_n1236_, new_n1237_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1256_, new_n1257_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1265_,
    new_n1266_, new_n1267_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1274_, new_n1275_, new_n1276_, new_n1278_, new_n1279_, new_n1281_,
    new_n1282_, new_n1283_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_;
  BUF_X1    g0000(.A(G141), .Z(G144));
  BUF_X1    g0001(.A(G293), .Z(G298));
  BUF_X1    g0002(.A(G3173), .Z(G973));
  INV_X1    g0003(.A(G545), .ZN(G594));
  INV_X1    g0004(.A(G348), .ZN(G599));
  INV_X1    g0005(.A(G366), .ZN(G600));
  INV_X1    g0006(.A(G552), .ZN(G849));
  INV_X1    g0007(.A(G562), .ZN(G850));
  NOR2_X1   g0008(.A1(G849), .A2(G850), .ZN(G601));
  INV_X1    g0009(.A(G549), .ZN(G602));
  INV_X1    g0010(.A(G545), .ZN(G603));
  INV_X1    g0011(.A(G545), .ZN(G604));
  XNOR2_X1  g0012(.A(KEYINPUT0), .B(G338), .ZN(G611));
  INV_X1    g0013(.A(G358), .ZN(G612));
  NAND2_X1  g0014(.A1(G141), .A2(G145), .ZN(new_n444_));
  XNOR2_X1  g0015(.A(new_n444_), .B(KEYINPUT1), .ZN(G810));
  INV_X1    g0016(.A(G245), .ZN(G848));
  INV_X1    g0017(.A(G559), .ZN(G851));
  AND2_X1   g0018(.A1(G1), .A2(G373), .ZN(G634));
  INV_X1    g0019(.A(G136), .ZN(new_n449_));
  NOR2_X1   g0020(.A1(new_n449_), .A2(G3173), .ZN(G815));
  INV_X1    g0021(.A(G2824), .ZN(new_n451_));
  NAND2_X1  g0022(.A1(new_n451_), .A2(G27), .ZN(G845));
  NAND2_X1  g0023(.A1(G386), .A2(G556), .ZN(G847));
  BUF_X1    g0024(.A(G137), .Z(G926));
  BUF_X1    g0025(.A(G141), .Z(G923));
  BUF_X1    g0026(.A(G1), .Z(G921));
  BUF_X1    g0027(.A(G549), .Z(G892));
  BUF_X1    g0028(.A(G299), .Z(G887));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G549), .Z(G606));
  NAND2_X1  g0030(.A1(G27), .A2(G31), .ZN(G809));
  INV_X1    g0031(.A(G809), .ZN(new_n461_));
  NAND2_X1  g0032(.A1(new_n461_), .A2(G140), .ZN(G656));
  XNOR2_X1  g0033(.A(KEYINPUT3), .B(G1), .ZN(G993));
  BUF_X1    g0034(.A(G1), .Z(G978));
  BUF_X1    g0035(.A(G1), .Z(G949));
  XNOR2_X1  g0036(.A(KEYINPUT4), .B(G1), .ZN(G939));
  BUF_X1    g0037(.A(G299), .Z(G889));
  INV_X1    g0038(.A(G299), .ZN(G593));
  OR2_X1    g0039(.A1(G86), .A2(G2358), .ZN(new_n469_));
  INV_X1    g0040(.A(G2358), .ZN(new_n470_));
  OAI211_X1 g0041(.A(new_n469_), .B(new_n461_), .C1(G87), .C2(new_n470_), .ZN(G636));
  OR2_X1    g0042(.A1(G88), .A2(G2358), .ZN(new_n472_));
  OAI211_X1 g0043(.A(new_n472_), .B(new_n461_), .C1(G34), .C2(new_n470_), .ZN(G704));
  OAI211_X1 g0044(.A(new_n472_), .B(new_n461_), .C1(G34), .C2(new_n470_), .ZN(G717));
  NAND2_X1  g0045(.A1(new_n461_), .A2(G83), .ZN(G820));
  INV_X1    g0046(.A(G141), .ZN(new_n476_));
  AOI21_X1  g0047(.A(G809), .B1(G24), .B2(new_n470_), .ZN(new_n477_));
  NAND2_X1  g0048(.A1(G25), .A2(G2358), .ZN(new_n478_));
  AOI21_X1  g0049(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(G639));
  AOI21_X1  g0050(.A(G809), .B1(G26), .B2(new_n470_), .ZN(new_n480_));
  NAND2_X1  g0051(.A1(G81), .A2(G2358), .ZN(new_n481_));
  AOI21_X1  g0052(.A(new_n476_), .B1(new_n480_), .B2(new_n481_), .ZN(G673));
  INV_X1    g0053(.A(G79), .ZN(new_n483_));
  OAI21_X1  g0054(.A(new_n461_), .B1(new_n483_), .B2(G2358), .ZN(new_n484_));
  INV_X1    g0055(.A(KEYINPUT5), .ZN(new_n485_));
  OR2_X1    g0056(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  AND2_X1   g0057(.A1(G23), .A2(G2358), .ZN(new_n487_));
  AOI22_X1  g0058(.A1(new_n484_), .A2(new_n485_), .B1(new_n461_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g0059(.A(new_n476_), .B1(new_n486_), .B2(new_n488_), .ZN(G707));
  AOI21_X1  g0060(.A(G809), .B1(G82), .B2(new_n470_), .ZN(new_n490_));
  NAND2_X1  g0061(.A1(G80), .A2(G2358), .ZN(new_n491_));
  AOI21_X1  g0062(.A(new_n476_), .B1(new_n490_), .B2(new_n491_), .ZN(G715));
  NAND2_X1  g0063(.A1(KEYINPUT6), .A2(G3552), .ZN(new_n493_));
  INV_X1    g0064(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g0065(.A1(KEYINPUT6), .A2(G3552), .ZN(new_n495_));
  NOR2_X1   g0066(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g0067(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g0068(.A1(new_n497_), .A2(G324), .A3(G503), .ZN(new_n498_));
  INV_X1    g0069(.A(G324), .ZN(new_n499_));
  INV_X1    g0070(.A(G3548), .ZN(new_n500_));
  AOI21_X1  g0071(.A(G503), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g0072(.A(new_n501_), .B1(new_n499_), .B2(G3546), .ZN(new_n502_));
  AND2_X1   g0073(.A1(new_n499_), .A2(G503), .ZN(new_n503_));
  INV_X1    g0074(.A(G3550), .ZN(new_n504_));
  AOI21_X1  g0075(.A(KEYINPUT8), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AND3_X1   g0076(.A1(new_n503_), .A2(KEYINPUT8), .A3(new_n504_), .ZN(new_n506_));
  OAI211_X1 g0077(.A(new_n498_), .B(new_n502_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g0078(.A(G341), .ZN(new_n508_));
  AOI21_X1  g0079(.A(G523), .B1(new_n508_), .B2(new_n500_), .ZN(new_n509_));
  OAI21_X1  g0080(.A(new_n509_), .B1(new_n508_), .B2(G3546), .ZN(new_n510_));
  NOR2_X1   g0081(.A1(new_n497_), .A2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g0082(.A(G523), .B1(new_n504_), .B2(G341), .ZN(new_n512_));
  OAI21_X1  g0083(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g0084(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g0085(.A(KEYINPUT7), .B(G351), .Z(new_n515_));
  INV_X1    g0086(.A(G351), .ZN(new_n516_));
  OAI22_X1  g0087(.A1(new_n515_), .A2(G3550), .B1(new_n496_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g0088(.A(G3546), .ZN(new_n518_));
  NAND2_X1  g0089(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g0090(.A(G534), .B1(new_n516_), .B2(new_n500_), .ZN(new_n520_));
  AOI22_X1  g0091(.A1(new_n517_), .A2(G534), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g0092(.A(G316), .ZN(new_n522_));
  AOI21_X1  g0093(.A(G490), .B1(new_n522_), .B2(G254), .ZN(new_n523_));
  INV_X1    g0094(.A(G242), .ZN(new_n524_));
  OAI21_X1  g0095(.A(new_n523_), .B1(new_n524_), .B2(new_n522_), .ZN(new_n525_));
  NOR2_X1   g0096(.A1(new_n522_), .A2(G248), .ZN(new_n526_));
  OAI21_X1  g0097(.A(G490), .B1(G251), .B2(G316), .ZN(new_n527_));
  OAI21_X1  g0098(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g0099(.A(G308), .ZN(new_n529_));
  AOI21_X1  g0100(.A(G479), .B1(new_n529_), .B2(G254), .ZN(new_n530_));
  OAI21_X1  g0101(.A(new_n530_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n531_));
  NOR2_X1   g0102(.A1(new_n529_), .A2(G248), .ZN(new_n532_));
  OAI21_X1  g0103(.A(G479), .B1(G251), .B2(G308), .ZN(new_n533_));
  OAI21_X1  g0104(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g0105(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g0106(.A1(G242), .A2(G293), .ZN(new_n536_));
  INV_X1    g0107(.A(G254), .ZN(new_n537_));
  OAI21_X1  g0108(.A(new_n536_), .B1(new_n537_), .B2(G293), .ZN(new_n538_));
  INV_X1    g0109(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g0110(.A(G514), .ZN(new_n540_));
  NAND2_X1  g0111(.A1(new_n540_), .A2(G3546), .ZN(new_n541_));
  OAI21_X1  g0112(.A(new_n541_), .B1(new_n540_), .B2(G3552), .ZN(new_n542_));
  NAND2_X1  g0113(.A1(G248), .A2(G302), .ZN(new_n543_));
  INV_X1    g0114(.A(G251), .ZN(new_n544_));
  OAI21_X1  g0115(.A(new_n543_), .B1(new_n544_), .B2(G302), .ZN(new_n545_));
  NAND2_X1  g0116(.A1(G248), .A2(G361), .ZN(new_n546_));
  OAI21_X1  g0117(.A(new_n546_), .B1(new_n544_), .B2(G361), .ZN(new_n547_));
  NAND4_X1  g0118(.A1(new_n539_), .A2(new_n542_), .A3(new_n545_), .A4(new_n547_), .ZN(new_n548_));
  NOR4_X1   g0119(.A1(new_n514_), .A2(new_n521_), .A3(new_n535_), .A4(new_n548_), .ZN(G598));
  INV_X1    g0120(.A(G281), .ZN(new_n550_));
  NOR2_X1   g0121(.A1(new_n497_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g0122(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g0123(.A(G374), .ZN(new_n553_));
  AOI21_X1  g0124(.A(new_n553_), .B1(new_n550_), .B2(G3550), .ZN(new_n554_));
  AOI21_X1  g0125(.A(G374), .B1(new_n518_), .B2(G281), .ZN(new_n555_));
  AOI22_X1  g0126(.A1(new_n555_), .A2(KEYINPUT13), .B1(new_n550_), .B2(new_n500_), .ZN(new_n556_));
  NOR2_X1   g0127(.A1(new_n555_), .A2(KEYINPUT13), .ZN(new_n557_));
  INV_X1    g0128(.A(new_n557_), .ZN(new_n558_));
  AOI22_X1  g0129(.A1(new_n552_), .A2(new_n554_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g0130(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g0131(.A(G389), .ZN(new_n561_));
  INV_X1    g0132(.A(G257), .ZN(new_n562_));
  AOI21_X1  g0133(.A(new_n561_), .B1(new_n562_), .B2(G3550), .ZN(new_n563_));
  OAI21_X1  g0134(.A(new_n563_), .B1(new_n497_), .B2(new_n562_), .ZN(new_n564_));
  OAI21_X1  g0135(.A(new_n561_), .B1(new_n562_), .B2(G3546), .ZN(new_n565_));
  AOI22_X1  g0136(.A1(new_n565_), .A2(KEYINPUT14), .B1(new_n562_), .B2(new_n500_), .ZN(new_n566_));
  OAI21_X1  g0137(.A(new_n566_), .B1(KEYINPUT14), .B2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g0138(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g0139(.A(G411), .ZN(new_n569_));
  INV_X1    g0140(.A(G273), .ZN(new_n570_));
  AOI21_X1  g0141(.A(new_n569_), .B1(new_n570_), .B2(G3550), .ZN(new_n571_));
  OAI21_X1  g0142(.A(new_n571_), .B1(new_n497_), .B2(new_n570_), .ZN(new_n572_));
  AOI21_X1  g0143(.A(G411), .B1(new_n570_), .B2(new_n500_), .ZN(new_n573_));
  OAI21_X1  g0144(.A(new_n573_), .B1(new_n570_), .B2(G3546), .ZN(new_n574_));
  NAND2_X1  g0145(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g0146(.A(G400), .ZN(new_n576_));
  INV_X1    g0147(.A(G265), .ZN(new_n577_));
  AOI21_X1  g0148(.A(new_n576_), .B1(new_n577_), .B2(G3550), .ZN(new_n578_));
  OAI21_X1  g0149(.A(new_n578_), .B1(new_n497_), .B2(new_n577_), .ZN(new_n579_));
  AOI21_X1  g0150(.A(G400), .B1(new_n577_), .B2(new_n500_), .ZN(new_n580_));
  OAI21_X1  g0151(.A(new_n580_), .B1(new_n577_), .B2(G3546), .ZN(new_n581_));
  NAND2_X1  g0152(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g0153(.A1(new_n560_), .A2(new_n568_), .A3(new_n575_), .A4(new_n582_), .ZN(new_n583_));
  OR2_X1    g0154(.A1(new_n583_), .A2(KEYINPUT15), .ZN(new_n584_));
  NAND3_X1  g0155(.A1(G206), .A2(G248), .A3(G446), .ZN(new_n585_));
  XOR2_X1   g0156(.A(new_n585_), .B(KEYINPUT16), .Z(new_n586_));
  INV_X1    g0157(.A(G446), .ZN(new_n587_));
  NOR3_X1   g0158(.A1(new_n544_), .A2(new_n587_), .A3(G206), .ZN(new_n588_));
  OAI21_X1  g0159(.A(new_n587_), .B1(new_n537_), .B2(G206), .ZN(new_n589_));
  AOI21_X1  g0160(.A(new_n589_), .B1(G206), .B2(G242), .ZN(new_n590_));
  OR3_X1    g0161(.A1(new_n586_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  XOR2_X1   g0162(.A(new_n591_), .B(KEYINPUT17), .Z(new_n592_));
  INV_X1    g0163(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g0164(.A(G435), .ZN(new_n594_));
  OR2_X1    g0165(.A1(new_n594_), .A2(G234), .ZN(new_n595_));
  OR2_X1    g0166(.A1(new_n595_), .A2(G3550), .ZN(new_n596_));
  NAND2_X1  g0167(.A1(G234), .A2(G435), .ZN(new_n597_));
  AOI21_X1  g0168(.A(G435), .B1(new_n518_), .B2(G234), .ZN(new_n598_));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n599_));
  OAI22_X1  g0170(.A1(new_n598_), .A2(new_n599_), .B1(G234), .B2(G3548), .ZN(new_n600_));
  AND2_X1   g0171(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  OAI221_X1 g0172(.A(new_n596_), .B1(new_n496_), .B2(new_n597_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  INV_X1    g0173(.A(G218), .ZN(new_n603_));
  AOI21_X1  g0174(.A(G468), .B1(new_n603_), .B2(new_n500_), .ZN(new_n604_));
  OAI21_X1  g0175(.A(new_n604_), .B1(new_n603_), .B2(G3546), .ZN(new_n605_));
  NAND2_X1  g0176(.A1(G218), .A2(G468), .ZN(new_n606_));
  INV_X1    g0177(.A(G468), .ZN(new_n607_));
  NOR2_X1   g0178(.A1(new_n607_), .A2(G218), .ZN(new_n608_));
  XNOR2_X1  g0179(.A(new_n608_), .B(KEYINPUT9), .ZN(new_n609_));
  OAI221_X1 g0180(.A(new_n605_), .B1(new_n496_), .B2(new_n606_), .C1(new_n609_), .C2(G3550), .ZN(new_n610_));
  INV_X1    g0181(.A(G226), .ZN(new_n611_));
  AOI21_X1  g0182(.A(G422), .B1(new_n611_), .B2(new_n500_), .ZN(new_n612_));
  OAI21_X1  g0183(.A(new_n612_), .B1(new_n611_), .B2(G3546), .ZN(new_n613_));
  NAND2_X1  g0184(.A1(new_n611_), .A2(G422), .ZN(new_n614_));
  NAND2_X1  g0185(.A1(G226), .A2(G422), .ZN(new_n615_));
  OAI221_X1 g0186(.A(new_n613_), .B1(G3550), .B2(new_n614_), .C1(new_n496_), .C2(new_n615_), .ZN(new_n616_));
  AND4_X1   g0187(.A1(new_n593_), .A2(new_n602_), .A3(new_n610_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g0188(.A1(new_n583_), .A2(KEYINPUT15), .ZN(new_n618_));
  INV_X1    g0189(.A(G457), .ZN(new_n619_));
  XNOR2_X1  g0190(.A(KEYINPUT11), .B(G210), .ZN(new_n620_));
  INV_X1    g0191(.A(new_n620_), .ZN(new_n621_));
  OAI221_X1 g0192(.A(new_n619_), .B1(G210), .B2(G3548), .C1(new_n621_), .C2(G3546), .ZN(new_n622_));
  INV_X1    g0193(.A(G210), .ZN(new_n623_));
  NOR2_X1   g0194(.A1(new_n496_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g0195(.A1(new_n620_), .A2(G3550), .ZN(new_n625_));
  OAI21_X1  g0196(.A(G457), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g0197(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g0198(.A(new_n627_), .B(KEYINPUT12), .ZN(new_n628_));
  AND4_X1   g0199(.A1(new_n584_), .A2(new_n617_), .A3(new_n618_), .A4(new_n628_), .ZN(G610));
  MUX2_X1   g0200(.A(G234), .B(G241), .S(G335), .Z(new_n630_));
  XOR2_X1   g0201(.A(new_n630_), .B(KEYINPUT21), .Z(new_n631_));
  XNOR2_X1  g0202(.A(new_n631_), .B(G435), .ZN(new_n632_));
  INV_X1    g0203(.A(G335), .ZN(new_n633_));
  NOR2_X1   g0204(.A1(new_n633_), .A2(G264), .ZN(new_n634_));
  NOR2_X1   g0205(.A1(G257), .A2(G335), .ZN(new_n635_));
  NOR3_X1   g0206(.A1(new_n634_), .A2(KEYINPUT18), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n637_));
  NAND2_X1  g0208(.A1(new_n562_), .A2(new_n633_), .ZN(new_n638_));
  INV_X1    g0209(.A(G264), .ZN(new_n639_));
  NAND2_X1  g0210(.A1(new_n639_), .A2(G335), .ZN(new_n640_));
  AOI21_X1  g0211(.A(new_n637_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g0212(.A(new_n561_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g0213(.A(KEYINPUT18), .B1(new_n634_), .B2(new_n635_), .ZN(new_n643_));
  NAND3_X1  g0214(.A1(new_n638_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n644_));
  NAND3_X1  g0215(.A1(new_n643_), .A2(new_n644_), .A3(G389), .ZN(new_n645_));
  NAND2_X1  g0216(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g0217(.A(new_n646_), .B(KEYINPUT19), .ZN(new_n647_));
  NAND2_X1  g0218(.A1(new_n632_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g0219(.A1(G288), .A2(G335), .ZN(new_n649_));
  INV_X1    g0220(.A(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g0221(.A(KEYINPUT20), .B(G335), .ZN(new_n651_));
  AOI21_X1  g0222(.A(new_n650_), .B1(new_n651_), .B2(G281), .ZN(new_n652_));
  INV_X1    g0223(.A(KEYINPUT23), .ZN(new_n653_));
  NOR2_X1   g0224(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI211_X1 g0225(.A(KEYINPUT23), .B(new_n650_), .C1(new_n651_), .C2(G281), .ZN(new_n655_));
  OAI21_X1  g0226(.A(G374), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  AND2_X1   g0227(.A1(KEYINPUT20), .A2(G335), .ZN(new_n657_));
  NOR2_X1   g0228(.A1(KEYINPUT20), .A2(G335), .ZN(new_n658_));
  NOR2_X1   g0229(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g0230(.A1(new_n659_), .A2(new_n550_), .ZN(new_n660_));
  OAI21_X1  g0231(.A(KEYINPUT23), .B1(new_n660_), .B2(new_n650_), .ZN(new_n661_));
  NAND2_X1  g0232(.A1(new_n652_), .A2(new_n653_), .ZN(new_n662_));
  NAND3_X1  g0233(.A1(new_n661_), .A2(new_n553_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g0234(.A1(G280), .A2(G335), .ZN(new_n664_));
  OAI211_X1 g0235(.A(new_n664_), .B(G411), .C1(new_n570_), .C2(G335), .ZN(new_n665_));
  INV_X1    g0236(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g0237(.A1(new_n633_), .A2(G273), .ZN(new_n667_));
  AOI21_X1  g0238(.A(G411), .B1(new_n667_), .B2(new_n664_), .ZN(new_n668_));
  OAI21_X1  g0239(.A(KEYINPUT22), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g0240(.A(new_n664_), .B1(new_n570_), .B2(G335), .ZN(new_n670_));
  NAND2_X1  g0241(.A1(new_n670_), .A2(new_n569_), .ZN(new_n671_));
  INV_X1    g0242(.A(KEYINPUT22), .ZN(new_n672_));
  NAND3_X1  g0243(.A1(new_n671_), .A2(new_n672_), .A3(new_n665_), .ZN(new_n673_));
  NAND2_X1  g0244(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g0245(.A1(new_n656_), .A2(new_n663_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g0246(.A1(new_n633_), .A2(G265), .ZN(new_n676_));
  NAND2_X1  g0247(.A1(G272), .A2(G335), .ZN(new_n677_));
  NAND2_X1  g0248(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g0249(.A1(new_n678_), .A2(G400), .ZN(new_n679_));
  INV_X1    g0250(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g0251(.A(G400), .B1(G272), .B2(G335), .ZN(new_n681_));
  INV_X1    g0252(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g0253(.A(new_n682_), .B1(new_n651_), .B2(G265), .ZN(new_n683_));
  NOR2_X1   g0254(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g0255(.A(new_n684_), .ZN(new_n685_));
  NOR3_X1   g0256(.A1(new_n648_), .A2(new_n675_), .A3(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g0257(.A(new_n686_), .B(KEYINPUT24), .ZN(new_n687_));
  INV_X1    g0258(.A(new_n687_), .ZN(new_n688_));
  AND2_X1   g0259(.A1(G233), .A2(G335), .ZN(new_n689_));
  AOI21_X1  g0260(.A(new_n689_), .B1(new_n651_), .B2(G226), .ZN(new_n690_));
  INV_X1    g0261(.A(G422), .ZN(new_n691_));
  OR2_X1    g0262(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g0263(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  AND2_X1   g0264(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g0265(.A(new_n694_), .B(KEYINPUT25), .ZN(new_n695_));
  NAND2_X1  g0266(.A1(G225), .A2(G335), .ZN(new_n696_));
  OAI21_X1  g0267(.A(new_n696_), .B1(new_n659_), .B2(new_n603_), .ZN(new_n697_));
  NAND2_X1  g0268(.A1(new_n697_), .A2(G468), .ZN(new_n698_));
  OAI211_X1 g0269(.A(new_n607_), .B(new_n696_), .C1(new_n659_), .C2(new_n603_), .ZN(new_n699_));
  NAND2_X1  g0270(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g0271(.A(new_n700_), .ZN(new_n701_));
  MUX2_X1   g0272(.A(G206), .B(G209), .S(G335), .Z(new_n702_));
  XOR2_X1   g0273(.A(new_n702_), .B(KEYINPUT26), .Z(new_n703_));
  XNOR2_X1  g0274(.A(new_n703_), .B(new_n587_), .ZN(new_n704_));
  NAND2_X1  g0275(.A1(new_n620_), .A2(new_n633_), .ZN(new_n705_));
  NAND2_X1  g0276(.A1(G217), .A2(G335), .ZN(new_n706_));
  NAND2_X1  g0277(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g0278(.A(new_n707_), .ZN(new_n708_));
  NOR2_X1   g0279(.A1(new_n708_), .A2(new_n619_), .ZN(new_n709_));
  NOR2_X1   g0280(.A1(new_n707_), .A2(G457), .ZN(new_n710_));
  NOR2_X1   g0281(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g0282(.A1(new_n695_), .A2(new_n701_), .A3(new_n704_), .A4(new_n711_), .ZN(new_n712_));
  NOR2_X1   g0283(.A1(new_n688_), .A2(new_n712_), .ZN(G588));
  MUX2_X1   g0284(.A(G324), .B(G331), .S(G332), .Z(new_n714_));
  XNOR2_X1  g0285(.A(new_n714_), .B(KEYINPUT30), .ZN(new_n715_));
  NOR2_X1   g0286(.A1(new_n715_), .A2(G503), .ZN(new_n716_));
  INV_X1    g0287(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g0288(.A1(new_n715_), .A2(G503), .ZN(new_n718_));
  AND2_X1   g0289(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g0290(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g0291(.A1(G611), .A2(G332), .ZN(new_n721_));
  NAND2_X1  g0292(.A1(new_n721_), .A2(KEYINPUT31), .ZN(new_n722_));
  INV_X1    g0293(.A(KEYINPUT31), .ZN(new_n723_));
  NAND3_X1  g0294(.A1(G611), .A2(new_n723_), .A3(G332), .ZN(new_n724_));
  NAND3_X1  g0295(.A1(new_n722_), .A2(new_n540_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g0296(.A1(new_n721_), .A2(G514), .ZN(new_n726_));
  NAND2_X1  g0297(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g0298(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g0299(.A1(G332), .A2(G348), .ZN(new_n729_));
  OAI21_X1  g0300(.A(new_n729_), .B1(new_n508_), .B2(G332), .ZN(new_n730_));
  INV_X1    g0301(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g0302(.A(G523), .ZN(new_n732_));
  NAND2_X1  g0303(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g0304(.A(new_n733_), .ZN(new_n734_));
  NOR2_X1   g0305(.A1(new_n731_), .A2(new_n732_), .ZN(new_n735_));
  NOR2_X1   g0306(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g0307(.A1(new_n728_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g0308(.A1(new_n720_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g0309(.A(G332), .ZN(new_n739_));
  NAND2_X1  g0310(.A1(new_n515_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g0311(.A1(G332), .A2(G358), .ZN(new_n741_));
  NAND2_X1  g0312(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g0313(.A(G534), .ZN(new_n743_));
  NAND2_X1  g0314(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g0315(.A1(new_n744_), .A2(KEYINPUT32), .ZN(new_n745_));
  OAI21_X1  g0316(.A(new_n741_), .B1(new_n516_), .B2(G332), .ZN(new_n746_));
  INV_X1    g0317(.A(new_n746_), .ZN(new_n747_));
  NAND2_X1  g0318(.A1(new_n747_), .A2(G534), .ZN(new_n748_));
  INV_X1    g0319(.A(KEYINPUT32), .ZN(new_n749_));
  NAND3_X1  g0320(.A1(new_n742_), .A2(new_n749_), .A3(new_n743_), .ZN(new_n750_));
  NAND3_X1  g0321(.A1(new_n745_), .A2(new_n748_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g0322(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g0323(.A1(G332), .A2(G366), .ZN(new_n753_));
  INV_X1    g0324(.A(G361), .ZN(new_n754_));
  OAI21_X1  g0325(.A(new_n753_), .B1(new_n754_), .B2(G332), .ZN(new_n755_));
  NOR2_X1   g0326(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g0327(.A1(new_n738_), .A2(new_n756_), .ZN(new_n757_));
  AND3_X1   g0328(.A1(KEYINPUT28), .A2(G315), .A3(G332), .ZN(new_n758_));
  OAI21_X1  g0329(.A(KEYINPUT28), .B1(new_n529_), .B2(G332), .ZN(new_n759_));
  NAND2_X1  g0330(.A1(G315), .A2(G332), .ZN(new_n760_));
  AOI21_X1  g0331(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g0332(.A(G479), .ZN(new_n762_));
  NAND2_X1  g0333(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g0334(.A(KEYINPUT29), .B(G479), .ZN(new_n764_));
  OAI21_X1  g0335(.A(new_n763_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g0336(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g0337(.A1(G323), .A2(G332), .ZN(new_n767_));
  OAI21_X1  g0338(.A(new_n767_), .B1(new_n522_), .B2(G332), .ZN(new_n768_));
  OR2_X1    g0339(.A1(new_n768_), .A2(G490), .ZN(new_n769_));
  NAND2_X1  g0340(.A1(new_n768_), .A2(G490), .ZN(new_n770_));
  NAND3_X1  g0341(.A1(new_n766_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g0342(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g0343(.A1(new_n739_), .A2(G302), .ZN(new_n773_));
  NAND2_X1  g0344(.A1(G307), .A2(G332), .ZN(new_n774_));
  AND2_X1   g0345(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g0346(.A1(G299), .A2(G332), .ZN(new_n776_));
  INV_X1    g0347(.A(G293), .ZN(new_n777_));
  OAI21_X1  g0348(.A(new_n776_), .B1(new_n777_), .B2(G332), .ZN(new_n778_));
  XNOR2_X1  g0349(.A(new_n778_), .B(KEYINPUT27), .ZN(new_n779_));
  NAND3_X1  g0350(.A1(new_n772_), .A2(new_n775_), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g0351(.A1(new_n757_), .A2(new_n780_), .ZN(G615));
  NOR2_X1   g0352(.A1(new_n757_), .A2(new_n780_), .ZN(G626));
  XNOR2_X1  g0353(.A(new_n631_), .B(new_n594_), .ZN(new_n783_));
  NAND2_X1  g0354(.A1(new_n656_), .A2(new_n663_), .ZN(new_n784_));
  INV_X1    g0355(.A(new_n784_), .ZN(new_n785_));
  AOI22_X1  g0356(.A1(new_n678_), .A2(G400), .B1(new_n676_), .B2(new_n681_), .ZN(new_n786_));
  NAND2_X1  g0357(.A1(new_n674_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g0358(.A1(new_n787_), .A2(new_n646_), .ZN(new_n788_));
  NAND2_X1  g0359(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NOR3_X1   g0360(.A1(new_n712_), .A2(new_n783_), .A3(new_n789_), .ZN(G632));
  XNOR2_X1  g0361(.A(G361), .B(G369), .ZN(new_n791_));
  XNOR2_X1  g0362(.A(new_n791_), .B(new_n499_), .ZN(new_n792_));
  XNOR2_X1  g0363(.A(G341), .B(G351), .ZN(new_n793_));
  XNOR2_X1  g0364(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g0365(.A(G293), .B(G302), .ZN(new_n795_));
  XNOR2_X1  g0366(.A(G308), .B(G316), .ZN(new_n796_));
  XNOR2_X1  g0367(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g0368(.A(new_n794_), .B(new_n797_), .ZN(G1002));
  XOR2_X1   g0369(.A(G206), .B(G210), .Z(new_n799_));
  XNOR2_X1  g0370(.A(KEYINPUT33), .B(G265), .ZN(new_n800_));
  XNOR2_X1  g0371(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g0372(.A(G218), .B(G226), .ZN(new_n802_));
  XNOR2_X1  g0373(.A(KEYINPUT34), .B(G273), .ZN(new_n803_));
  XNOR2_X1  g0374(.A(new_n802_), .B(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g0375(.A(new_n801_), .B(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g0376(.A(G234), .B(G257), .ZN(new_n806_));
  XNOR2_X1  g0377(.A(G281), .B(G289), .ZN(new_n807_));
  XNOR2_X1  g0378(.A(new_n806_), .B(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g0379(.A(new_n805_), .B(new_n808_), .ZN(G1004));
  NAND2_X1  g0380(.A1(new_n703_), .A2(G446), .ZN(new_n810_));
  INV_X1    g0381(.A(new_n704_), .ZN(new_n811_));
  NOR2_X1   g0382(.A1(new_n690_), .A2(new_n691_), .ZN(new_n812_));
  NAND2_X1  g0383(.A1(new_n812_), .A2(new_n699_), .ZN(new_n813_));
  NAND2_X1  g0384(.A1(new_n813_), .A2(new_n698_), .ZN(new_n814_));
  INV_X1    g0385(.A(new_n710_), .ZN(new_n815_));
  AOI21_X1  g0386(.A(new_n709_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OR2_X1    g0387(.A1(new_n631_), .A2(new_n594_), .ZN(new_n817_));
  XNOR2_X1  g0388(.A(new_n645_), .B(KEYINPUT35), .ZN(new_n818_));
  AOI21_X1  g0389(.A(new_n818_), .B1(new_n594_), .B2(new_n631_), .ZN(new_n819_));
  NAND2_X1  g0390(.A1(new_n651_), .A2(G281), .ZN(new_n820_));
  AOI21_X1  g0391(.A(new_n553_), .B1(new_n820_), .B2(new_n649_), .ZN(new_n821_));
  NOR3_X1   g0392(.A1(new_n666_), .A2(new_n668_), .A3(KEYINPUT22), .ZN(new_n822_));
  AOI21_X1  g0393(.A(new_n672_), .B1(new_n671_), .B2(new_n665_), .ZN(new_n823_));
  OAI211_X1 g0394(.A(new_n786_), .B(new_n821_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n824_));
  OAI221_X1 g0395(.A(new_n817_), .B1(new_n819_), .B2(KEYINPUT36), .C1(new_n648_), .C2(new_n824_), .ZN(new_n825_));
  XOR2_X1   g0396(.A(new_n645_), .B(KEYINPUT35), .Z(new_n826_));
  NAND2_X1  g0397(.A1(new_n826_), .A2(KEYINPUT36), .ZN(new_n827_));
  AND2_X1   g0398(.A1(new_n642_), .A2(new_n645_), .ZN(new_n828_));
  OAI21_X1  g0399(.A(G273), .B1(new_n657_), .B2(new_n658_), .ZN(new_n829_));
  AOI21_X1  g0400(.A(new_n569_), .B1(new_n829_), .B2(new_n664_), .ZN(new_n830_));
  AND2_X1   g0401(.A1(new_n830_), .A2(new_n786_), .ZN(new_n831_));
  OAI21_X1  g0402(.A(new_n828_), .B1(new_n680_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g0403(.A(new_n783_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g0404(.A1(new_n825_), .A2(new_n833_), .ZN(new_n834_));
  OAI221_X1 g0405(.A(new_n810_), .B1(new_n811_), .B2(new_n816_), .C1(new_n834_), .C2(new_n712_), .ZN(G591));
  NOR2_X1   g0406(.A1(new_n761_), .A2(new_n762_), .ZN(new_n836_));
  XNOR2_X1  g0407(.A(new_n770_), .B(KEYINPUT37), .ZN(new_n837_));
  AOI21_X1  g0408(.A(new_n836_), .B1(new_n766_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g0409(.A1(new_n838_), .A2(new_n775_), .ZN(new_n839_));
  NOR2_X1   g0410(.A1(new_n839_), .A2(new_n778_), .ZN(new_n840_));
  AOI21_X1  g0411(.A(new_n540_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n841_));
  NAND3_X1  g0412(.A1(new_n745_), .A2(new_n743_), .A3(new_n750_), .ZN(new_n842_));
  INV_X1    g0413(.A(new_n755_), .ZN(new_n843_));
  OAI21_X1  g0414(.A(new_n843_), .B1(new_n747_), .B2(new_n743_), .ZN(new_n844_));
  NAND3_X1  g0415(.A1(new_n842_), .A2(new_n733_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g0416(.A(new_n735_), .ZN(new_n846_));
  NAND2_X1  g0417(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g0418(.A(new_n841_), .B1(new_n847_), .B2(new_n728_), .ZN(new_n848_));
  OAI21_X1  g0419(.A(new_n718_), .B1(new_n848_), .B2(new_n716_), .ZN(new_n849_));
  XNOR2_X1  g0420(.A(new_n849_), .B(KEYINPUT38), .ZN(new_n850_));
  OAI21_X1  g0421(.A(new_n840_), .B1(new_n850_), .B2(new_n780_), .ZN(G618));
  OAI221_X1 g0422(.A(new_n810_), .B1(new_n811_), .B2(new_n816_), .C1(new_n834_), .C2(new_n712_), .ZN(G621));
  OAI21_X1  g0423(.A(new_n840_), .B1(new_n850_), .B2(new_n780_), .ZN(G629));
  INV_X1    g0424(.A(G4092), .ZN(new_n854_));
  NOR2_X1   g0425(.A1(new_n854_), .A2(G4091), .ZN(new_n855_));
  NAND2_X1  g0426(.A1(new_n855_), .A2(G131), .ZN(new_n856_));
  NOR2_X1   g0427(.A1(G4091), .A2(G4092), .ZN(new_n857_));
  INV_X1    g0428(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g0429(.A(G54), .ZN(new_n859_));
  XNOR2_X1  g0430(.A(new_n755_), .B(new_n859_), .ZN(new_n860_));
  INV_X1    g0431(.A(G4091), .ZN(new_n861_));
  NOR2_X1   g0432(.A1(new_n861_), .A2(G4092), .ZN(new_n862_));
  INV_X1    g0433(.A(new_n862_), .ZN(new_n863_));
  OAI221_X1 g0434(.A(new_n856_), .B1(new_n547_), .B2(new_n858_), .C1(new_n860_), .C2(new_n863_), .ZN(new_n864_));
  INV_X1    g0435(.A(new_n864_), .ZN(G822));
  AOI22_X1  g0436(.A1(new_n521_), .A2(new_n857_), .B1(G129), .B2(new_n855_), .ZN(new_n866_));
  NAND2_X1  g0437(.A1(new_n843_), .A2(new_n859_), .ZN(new_n867_));
  INV_X1    g0438(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g0439(.A(new_n863_), .B1(new_n752_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g0440(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g0441(.A1(new_n752_), .A2(new_n868_), .ZN(new_n871_));
  OAI21_X1  g0442(.A(new_n866_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g0443(.A(new_n872_), .ZN(G838));
  XNOR2_X1  g0444(.A(new_n784_), .B(G4), .ZN(new_n874_));
  NAND2_X1  g0445(.A1(new_n874_), .A2(new_n862_), .ZN(new_n875_));
  NAND2_X1  g0446(.A1(new_n560_), .A2(new_n854_), .ZN(new_n876_));
  OAI211_X1 g0447(.A(new_n876_), .B(new_n861_), .C1(G117), .C2(new_n854_), .ZN(new_n877_));
  NAND2_X1  g0448(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g0449(.A(new_n878_), .ZN(G861));
  NAND3_X1  g0450(.A1(new_n738_), .A2(G54), .A3(new_n756_), .ZN(new_n880_));
  NAND2_X1  g0451(.A1(new_n850_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g0452(.A(KEYINPUT39), .ZN(new_n882_));
  NAND2_X1  g0453(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g0454(.A1(new_n850_), .A2(KEYINPUT39), .A3(new_n880_), .ZN(new_n884_));
  NAND2_X1  g0455(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g0456(.A(new_n769_), .ZN(new_n886_));
  OAI221_X1 g0457(.A(new_n775_), .B1(new_n762_), .B2(new_n761_), .C1(new_n765_), .C2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g0458(.A(new_n887_), .B(new_n778_), .ZN(new_n888_));
  NAND2_X1  g0459(.A1(new_n885_), .A2(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g0460(.A(new_n839_), .B(KEYINPUT40), .ZN(new_n890_));
  XOR2_X1   g0461(.A(new_n890_), .B(new_n779_), .Z(new_n891_));
  OAI21_X1  g0462(.A(new_n889_), .B1(new_n885_), .B2(new_n891_), .ZN(new_n892_));
  XOR2_X1   g0463(.A(new_n892_), .B(KEYINPUT41), .Z(new_n893_));
  INV_X1    g0464(.A(new_n893_), .ZN(G623));
  OAI21_X1  g0465(.A(G4087), .B1(G11), .B2(G4088), .ZN(new_n895_));
  INV_X1    g0466(.A(G61), .ZN(new_n896_));
  AOI21_X1  g0467(.A(new_n895_), .B1(new_n896_), .B2(G4088), .ZN(new_n897_));
  NOR2_X1   g0468(.A1(G4087), .A2(G4088), .ZN(new_n898_));
  AOI21_X1  g0469(.A(new_n897_), .B1(new_n864_), .B2(new_n898_), .ZN(new_n899_));
  XOR2_X1   g0470(.A(new_n878_), .B(KEYINPUT42), .Z(new_n900_));
  XNOR2_X1  g0471(.A(KEYINPUT43), .B(G4087), .ZN(new_n901_));
  INV_X1    g0472(.A(G4088), .ZN(new_n902_));
  NOR2_X1   g0473(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g0474(.A(new_n903_), .ZN(new_n904_));
  OAI21_X1  g0475(.A(new_n899_), .B1(new_n900_), .B2(new_n904_), .ZN(G722));
  NAND2_X1  g0476(.A1(new_n507_), .A2(new_n854_), .ZN(new_n906_));
  OAI211_X1 g0477(.A(new_n906_), .B(new_n861_), .C1(G52), .C2(new_n854_), .ZN(new_n907_));
  NAND4_X1  g0478(.A1(new_n751_), .A2(new_n736_), .A3(new_n728_), .A4(new_n755_), .ZN(new_n908_));
  NAND3_X1  g0479(.A1(new_n733_), .A2(G534), .A3(new_n746_), .ZN(new_n909_));
  NAND2_X1  g0480(.A1(new_n909_), .A2(new_n846_), .ZN(new_n910_));
  AOI21_X1  g0481(.A(new_n841_), .B1(new_n728_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g0482(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g0483(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g0484(.A1(new_n756_), .A2(G54), .ZN(new_n914_));
  OAI21_X1  g0485(.A(new_n913_), .B1(new_n914_), .B2(new_n737_), .ZN(new_n915_));
  XNOR2_X1  g0486(.A(new_n915_), .B(new_n719_), .ZN(new_n916_));
  OAI21_X1  g0487(.A(new_n907_), .B1(new_n916_), .B2(new_n863_), .ZN(new_n917_));
  XNOR2_X1  g0488(.A(new_n917_), .B(KEYINPUT44), .ZN(new_n918_));
  INV_X1    g0489(.A(new_n918_), .ZN(G832));
  OAI21_X1  g0490(.A(new_n861_), .B1(new_n854_), .B2(G130), .ZN(new_n920_));
  AOI21_X1  g0491(.A(new_n920_), .B1(new_n542_), .B2(new_n854_), .ZN(new_n921_));
  AOI21_X1  g0492(.A(new_n910_), .B1(new_n871_), .B2(new_n733_), .ZN(new_n922_));
  XNOR2_X1  g0493(.A(new_n922_), .B(new_n728_), .ZN(new_n923_));
  AOI21_X1  g0494(.A(new_n921_), .B1(new_n923_), .B2(new_n862_), .ZN(G834));
  NAND2_X1  g0495(.A1(new_n747_), .A2(new_n743_), .ZN(new_n925_));
  NAND2_X1  g0496(.A1(new_n844_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g0497(.A1(new_n914_), .A2(new_n926_), .ZN(new_n927_));
  XOR2_X1   g0498(.A(new_n736_), .B(KEYINPUT45), .Z(new_n928_));
  XNOR2_X1  g0499(.A(new_n927_), .B(new_n928_), .ZN(new_n929_));
  NOR2_X1   g0500(.A1(new_n929_), .A2(new_n863_), .ZN(new_n930_));
  OAI21_X1  g0501(.A(new_n861_), .B1(new_n854_), .B2(G119), .ZN(new_n931_));
  AOI21_X1  g0502(.A(new_n931_), .B1(new_n513_), .B2(new_n854_), .ZN(new_n932_));
  NOR2_X1   g0503(.A1(new_n930_), .A2(new_n932_), .ZN(G836));
  OAI21_X1  g0504(.A(G4090), .B1(G11), .B2(G4089), .ZN(new_n934_));
  AOI21_X1  g0505(.A(new_n934_), .B1(new_n896_), .B2(G4089), .ZN(new_n935_));
  NOR2_X1   g0506(.A1(G4089), .A2(G4090), .ZN(new_n936_));
  AOI21_X1  g0507(.A(new_n935_), .B1(new_n864_), .B2(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g0508(.A(KEYINPUT46), .B(G4090), .ZN(new_n938_));
  INV_X1    g0509(.A(G4089), .ZN(new_n939_));
  NOR2_X1   g0510(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g0511(.A(new_n940_), .ZN(new_n941_));
  OAI21_X1  g0512(.A(new_n937_), .B1(new_n900_), .B2(new_n941_), .ZN(G859));
  NOR2_X1   g0513(.A1(new_n646_), .A2(new_n679_), .ZN(new_n943_));
  NAND4_X1  g0514(.A1(new_n831_), .A2(KEYINPUT47), .A3(new_n645_), .A4(new_n642_), .ZN(new_n944_));
  INV_X1    g0515(.A(KEYINPUT47), .ZN(new_n945_));
  NAND2_X1  g0516(.A1(new_n830_), .A2(new_n786_), .ZN(new_n946_));
  OAI21_X1  g0517(.A(new_n945_), .B1(new_n646_), .B2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g0518(.A1(new_n944_), .A2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g0519(.A1(new_n681_), .A2(new_n676_), .ZN(new_n949_));
  NAND2_X1  g0520(.A1(new_n679_), .A2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g0521(.A(new_n950_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n951_));
  INV_X1    g0522(.A(KEYINPUT48), .ZN(new_n952_));
  NAND4_X1  g0523(.A1(new_n828_), .A2(new_n951_), .A3(new_n952_), .A4(new_n821_), .ZN(new_n953_));
  OAI21_X1  g0524(.A(KEYINPUT48), .B1(new_n824_), .B2(new_n646_), .ZN(new_n954_));
  AOI21_X1  g0525(.A(new_n948_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g0526(.A(G4), .ZN(new_n956_));
  NOR2_X1   g0527(.A1(new_n784_), .A2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g0528(.A1(new_n957_), .A2(new_n788_), .ZN(new_n958_));
  NAND2_X1  g0529(.A1(new_n955_), .A2(new_n958_), .ZN(new_n959_));
  AOI211_X1 g0530(.A(new_n826_), .B(new_n943_), .C1(new_n959_), .C2(KEYINPUT49), .ZN(new_n960_));
  OAI21_X1  g0531(.A(new_n960_), .B1(KEYINPUT49), .B2(new_n959_), .ZN(new_n961_));
  XNOR2_X1  g0532(.A(new_n961_), .B(new_n783_), .ZN(new_n962_));
  AND2_X1   g0533(.A1(new_n962_), .A2(new_n862_), .ZN(new_n963_));
  OAI21_X1  g0534(.A(new_n861_), .B1(new_n854_), .B2(G122), .ZN(new_n964_));
  AOI21_X1  g0535(.A(new_n964_), .B1(new_n602_), .B2(new_n854_), .ZN(new_n965_));
  NOR2_X1   g0536(.A1(new_n963_), .A2(new_n965_), .ZN(G871));
  NAND2_X1  g0537(.A1(new_n957_), .A2(new_n951_), .ZN(new_n967_));
  INV_X1    g0538(.A(KEYINPUT50), .ZN(new_n968_));
  NAND3_X1  g0539(.A1(new_n951_), .A2(new_n968_), .A3(new_n821_), .ZN(new_n969_));
  INV_X1    g0540(.A(new_n830_), .ZN(new_n970_));
  OAI21_X1  g0541(.A(new_n679_), .B1(new_n970_), .B2(new_n683_), .ZN(new_n971_));
  INV_X1    g0542(.A(new_n971_), .ZN(new_n972_));
  NAND2_X1  g0543(.A1(new_n824_), .A2(KEYINPUT50), .ZN(new_n973_));
  NAND4_X1  g0544(.A1(new_n967_), .A2(new_n969_), .A3(new_n972_), .A4(new_n973_), .ZN(new_n974_));
  XNOR2_X1  g0545(.A(new_n974_), .B(new_n828_), .ZN(new_n975_));
  OR2_X1    g0546(.A1(new_n975_), .A2(new_n863_), .ZN(new_n976_));
  NOR2_X1   g0547(.A1(new_n568_), .A2(G4092), .ZN(new_n977_));
  AND2_X1   g0548(.A1(new_n977_), .A2(KEYINPUT51), .ZN(new_n978_));
  NAND2_X1  g0549(.A1(G128), .A2(G4092), .ZN(new_n979_));
  OAI21_X1  g0550(.A(new_n979_), .B1(new_n977_), .B2(KEYINPUT51), .ZN(new_n980_));
  OAI21_X1  g0551(.A(new_n861_), .B1(new_n978_), .B2(new_n980_), .ZN(new_n981_));
  NAND2_X1  g0552(.A1(new_n976_), .A2(new_n981_), .ZN(new_n982_));
  INV_X1    g0553(.A(new_n982_), .ZN(G873));
  NAND2_X1  g0554(.A1(new_n829_), .A2(new_n664_), .ZN(new_n984_));
  NAND2_X1  g0555(.A1(new_n984_), .A2(new_n569_), .ZN(new_n985_));
  NAND2_X1  g0556(.A1(new_n985_), .A2(new_n665_), .ZN(new_n986_));
  NAND2_X1  g0557(.A1(new_n986_), .A2(new_n821_), .ZN(new_n987_));
  OR2_X1    g0558(.A1(new_n830_), .A2(KEYINPUT52), .ZN(new_n988_));
  NAND2_X1  g0559(.A1(new_n830_), .A2(KEYINPUT52), .ZN(new_n989_));
  NAND3_X1  g0560(.A1(new_n987_), .A2(new_n988_), .A3(new_n989_), .ZN(new_n990_));
  AOI21_X1  g0561(.A(new_n990_), .B1(new_n957_), .B2(new_n674_), .ZN(new_n991_));
  XNOR2_X1  g0562(.A(new_n786_), .B(KEYINPUT53), .ZN(new_n992_));
  XNOR2_X1  g0563(.A(new_n991_), .B(new_n992_), .ZN(new_n993_));
  NOR2_X1   g0564(.A1(new_n993_), .A2(new_n863_), .ZN(new_n994_));
  OAI21_X1  g0565(.A(new_n861_), .B1(new_n854_), .B2(G127), .ZN(new_n995_));
  AOI21_X1  g0566(.A(new_n995_), .B1(new_n582_), .B2(new_n854_), .ZN(new_n996_));
  NOR2_X1   g0567(.A1(new_n994_), .A2(new_n996_), .ZN(G875));
  NOR2_X1   g0568(.A1(new_n957_), .A2(new_n821_), .ZN(new_n998_));
  XNOR2_X1  g0569(.A(new_n998_), .B(new_n674_), .ZN(new_n999_));
  AND2_X1   g0570(.A1(new_n999_), .A2(new_n862_), .ZN(new_n1000_));
  NAND3_X1  g0571(.A1(new_n572_), .A2(new_n854_), .A3(new_n574_), .ZN(new_n1001_));
  OR2_X1    g0572(.A1(new_n1001_), .A2(KEYINPUT54), .ZN(new_n1002_));
  AOI22_X1  g0573(.A1(new_n1001_), .A2(KEYINPUT54), .B1(G126), .B2(G4092), .ZN(new_n1003_));
  AOI21_X1  g0574(.A(G4091), .B1(new_n1002_), .B2(new_n1003_), .ZN(new_n1004_));
  NOR2_X1   g0575(.A1(new_n1000_), .A2(new_n1004_), .ZN(G877));
  XNOR2_X1  g0576(.A(new_n715_), .B(new_n742_), .ZN(new_n1006_));
  MUX2_X1   g0577(.A(G369), .B(G372), .S(G332), .Z(new_n1007_));
  XNOR2_X1  g0578(.A(new_n1006_), .B(new_n1007_), .ZN(new_n1008_));
  XNOR2_X1  g0579(.A(new_n1008_), .B(new_n761_), .ZN(new_n1009_));
  NAND2_X1  g0580(.A1(new_n722_), .A2(new_n724_), .ZN(new_n1010_));
  XNOR2_X1  g0581(.A(new_n1010_), .B(new_n775_), .ZN(new_n1011_));
  XOR2_X1   g0582(.A(new_n768_), .B(new_n778_), .Z(new_n1012_));
  XNOR2_X1  g0583(.A(new_n1011_), .B(new_n1012_), .ZN(new_n1013_));
  XOR2_X1   g0584(.A(new_n755_), .B(KEYINPUT56), .Z(new_n1014_));
  XNOR2_X1  g0585(.A(new_n730_), .B(KEYINPUT55), .ZN(new_n1015_));
  XNOR2_X1  g0586(.A(new_n1014_), .B(new_n1015_), .ZN(new_n1016_));
  XNOR2_X1  g0587(.A(new_n1013_), .B(new_n1016_), .ZN(new_n1017_));
  XNOR2_X1  g0588(.A(new_n1009_), .B(new_n1017_), .ZN(G998));
  NAND2_X1  g0589(.A1(new_n661_), .A2(new_n662_), .ZN(new_n1019_));
  XNOR2_X1  g0590(.A(new_n1019_), .B(new_n708_), .ZN(new_n1020_));
  XNOR2_X1  g0591(.A(new_n678_), .B(new_n670_), .ZN(new_n1021_));
  XNOR2_X1  g0592(.A(new_n1020_), .B(new_n1021_), .ZN(new_n1022_));
  MUX2_X1   g0593(.A(G289), .B(G292), .S(G335), .Z(new_n1023_));
  XNOR2_X1  g0594(.A(new_n631_), .B(new_n1023_), .ZN(new_n1024_));
  XNOR2_X1  g0595(.A(new_n1022_), .B(new_n1024_), .ZN(new_n1025_));
  XNOR2_X1  g0596(.A(new_n703_), .B(KEYINPUT57), .ZN(new_n1026_));
  XNOR2_X1  g0597(.A(new_n1026_), .B(new_n690_), .ZN(new_n1027_));
  XNOR2_X1  g0598(.A(new_n697_), .B(KEYINPUT58), .ZN(new_n1028_));
  NAND2_X1  g0599(.A1(new_n643_), .A2(new_n644_), .ZN(new_n1029_));
  XOR2_X1   g0600(.A(new_n1028_), .B(new_n1029_), .Z(new_n1030_));
  XNOR2_X1  g0601(.A(new_n1027_), .B(new_n1030_), .ZN(new_n1031_));
  XNOR2_X1  g0602(.A(new_n1025_), .B(new_n1031_), .ZN(G1000));
  NOR2_X1   g0603(.A1(new_n789_), .A2(new_n783_), .ZN(new_n1033_));
  AOI21_X1  g0604(.A(new_n956_), .B1(new_n1033_), .B2(KEYINPUT59), .ZN(new_n1034_));
  OAI21_X1  g0605(.A(new_n1034_), .B1(KEYINPUT59), .B2(new_n1033_), .ZN(new_n1035_));
  NAND2_X1  g0606(.A1(new_n1035_), .A2(new_n834_), .ZN(new_n1036_));
  XNOR2_X1  g0607(.A(new_n1036_), .B(KEYINPUT60), .ZN(new_n1037_));
  XNOR2_X1  g0608(.A(new_n1037_), .B(KEYINPUT61), .ZN(new_n1038_));
  INV_X1    g0609(.A(new_n1038_), .ZN(new_n1039_));
  XNOR2_X1  g0610(.A(new_n816_), .B(new_n704_), .ZN(new_n1040_));
  INV_X1    g0611(.A(new_n1037_), .ZN(new_n1041_));
  INV_X1    g0612(.A(new_n709_), .ZN(new_n1042_));
  NAND2_X1  g0613(.A1(new_n693_), .A2(new_n699_), .ZN(new_n1043_));
  AND2_X1   g0614(.A1(new_n1043_), .A2(new_n698_), .ZN(new_n1044_));
  OAI21_X1  g0615(.A(new_n1042_), .B1(new_n1044_), .B2(new_n710_), .ZN(new_n1045_));
  XNOR2_X1  g0616(.A(new_n811_), .B(new_n1045_), .ZN(new_n1046_));
  AOI22_X1  g0617(.A1(new_n1039_), .A2(new_n1040_), .B1(new_n1041_), .B2(new_n1046_), .ZN(new_n1047_));
  INV_X1    g0618(.A(new_n695_), .ZN(new_n1048_));
  XNOR2_X1  g0619(.A(new_n1037_), .B(new_n1048_), .ZN(new_n1049_));
  NAND2_X1  g0620(.A1(new_n1047_), .A2(new_n1049_), .ZN(new_n1050_));
  XOR2_X1   g0621(.A(new_n711_), .B(new_n814_), .Z(new_n1051_));
  NAND2_X1  g0622(.A1(new_n1039_), .A2(new_n1051_), .ZN(new_n1052_));
  XNOR2_X1  g0623(.A(new_n711_), .B(new_n1044_), .ZN(new_n1053_));
  NAND2_X1  g0624(.A1(new_n1041_), .A2(new_n1053_), .ZN(new_n1054_));
  NAND2_X1  g0625(.A1(new_n1052_), .A2(new_n1054_), .ZN(new_n1055_));
  AOI21_X1  g0626(.A(new_n1050_), .B1(KEYINPUT62), .B2(new_n1055_), .ZN(new_n1056_));
  OAI21_X1  g0627(.A(new_n693_), .B1(new_n1038_), .B2(new_n812_), .ZN(new_n1057_));
  XNOR2_X1  g0628(.A(new_n1057_), .B(new_n701_), .ZN(new_n1058_));
  INV_X1    g0629(.A(new_n1058_), .ZN(new_n1059_));
  OAI211_X1 g0630(.A(new_n1056_), .B(new_n1059_), .C1(KEYINPUT62), .C2(new_n1055_), .ZN(new_n1060_));
  XNOR2_X1  g0631(.A(new_n1060_), .B(KEYINPUT63), .ZN(new_n1061_));
  NOR2_X1   g0632(.A1(new_n999_), .A2(new_n874_), .ZN(new_n1062_));
  NAND3_X1  g0633(.A1(new_n975_), .A2(new_n1062_), .A3(new_n993_), .ZN(new_n1063_));
  NOR3_X1   g0634(.A1(new_n1061_), .A2(new_n962_), .A3(new_n1063_), .ZN(G575));
  INV_X1    g0635(.A(new_n885_), .ZN(new_n1065_));
  NAND2_X1  g0636(.A1(new_n1065_), .A2(new_n837_), .ZN(new_n1066_));
  OAI21_X1  g0637(.A(new_n1066_), .B1(new_n886_), .B2(new_n1065_), .ZN(new_n1067_));
  XNOR2_X1  g0638(.A(new_n1067_), .B(new_n765_), .ZN(new_n1068_));
  NAND2_X1  g0639(.A1(new_n769_), .A2(new_n770_), .ZN(new_n1069_));
  XOR2_X1   g0640(.A(new_n885_), .B(new_n1069_), .Z(new_n1070_));
  INV_X1    g0641(.A(new_n1070_), .ZN(new_n1071_));
  OAI21_X1  g0642(.A(new_n838_), .B1(new_n1065_), .B2(new_n771_), .ZN(new_n1072_));
  INV_X1    g0643(.A(new_n775_), .ZN(new_n1073_));
  XNOR2_X1  g0644(.A(new_n1072_), .B(new_n1073_), .ZN(new_n1074_));
  NOR4_X1   g0645(.A1(new_n1068_), .A2(new_n893_), .A3(new_n1071_), .A4(new_n1074_), .ZN(new_n1075_));
  XNOR2_X1  g0646(.A(new_n1075_), .B(KEYINPUT64), .ZN(new_n1076_));
  INV_X1    g0647(.A(new_n860_), .ZN(new_n1077_));
  NOR3_X1   g0648(.A1(new_n923_), .A2(new_n752_), .A3(new_n1077_), .ZN(new_n1078_));
  AND4_X1   g0649(.A1(new_n916_), .A2(new_n1076_), .A3(new_n929_), .A4(new_n1078_), .ZN(G585));
  INV_X1    g0650(.A(G137), .ZN(new_n1080_));
  INV_X1    g0651(.A(G1689), .ZN(new_n1081_));
  NOR2_X1   g0652(.A1(new_n1081_), .A2(G1690), .ZN(new_n1082_));
  INV_X1    g0653(.A(new_n1082_), .ZN(new_n1083_));
  NOR2_X1   g0654(.A1(new_n900_), .A2(new_n1083_), .ZN(new_n1084_));
  XNOR2_X1  g0655(.A(new_n1084_), .B(KEYINPUT65), .ZN(new_n1085_));
  OAI21_X1  g0656(.A(G1690), .B1(G182), .B2(G1689), .ZN(new_n1086_));
  INV_X1    g0657(.A(G185), .ZN(new_n1087_));
  AOI21_X1  g0658(.A(new_n1086_), .B1(new_n1087_), .B2(G1689), .ZN(new_n1088_));
  NOR2_X1   g0659(.A1(G1689), .A2(G1690), .ZN(new_n1089_));
  AOI21_X1  g0660(.A(new_n1088_), .B1(new_n864_), .B2(new_n1089_), .ZN(new_n1090_));
  AOI21_X1  g0661(.A(new_n1080_), .B1(new_n1085_), .B2(new_n1090_), .ZN(G661));
  INV_X1    g0662(.A(G1694), .ZN(new_n1092_));
  NAND2_X1  g0663(.A1(new_n864_), .A2(new_n1092_), .ZN(new_n1093_));
  OAI21_X1  g0664(.A(G1694), .B1(G182), .B2(G1691), .ZN(new_n1094_));
  AND3_X1   g0665(.A1(new_n1093_), .A2(KEYINPUT66), .A3(new_n1094_), .ZN(new_n1095_));
  INV_X1    g0666(.A(G1691), .ZN(new_n1096_));
  OAI21_X1  g0667(.A(new_n1096_), .B1(new_n1093_), .B2(KEYINPUT66), .ZN(new_n1097_));
  OAI22_X1  g0668(.A1(new_n1095_), .A2(new_n1097_), .B1(new_n1087_), .B2(new_n1094_), .ZN(new_n1098_));
  INV_X1    g0669(.A(new_n900_), .ZN(new_n1099_));
  NOR2_X1   g0670(.A1(new_n1096_), .A2(G1694), .ZN(new_n1100_));
  AOI21_X1  g0671(.A(new_n1098_), .B1(new_n1099_), .B2(new_n1100_), .ZN(new_n1101_));
  NOR2_X1   g0672(.A1(new_n1101_), .A2(new_n1080_), .ZN(new_n1102_));
  XNOR2_X1  g0673(.A(new_n1102_), .B(KEYINPUT67), .ZN(G693));
  OR2_X1    g0674(.A1(G43), .A2(G4088), .ZN(new_n1104_));
  OAI211_X1 g0675(.A(new_n1104_), .B(G4087), .C1(G37), .C2(new_n902_), .ZN(new_n1105_));
  NOR2_X1   g0676(.A1(new_n901_), .A2(G4088), .ZN(new_n1106_));
  INV_X1    g0677(.A(new_n1106_), .ZN(new_n1107_));
  OAI221_X1 g0678(.A(new_n1105_), .B1(G832), .B2(new_n1107_), .C1(new_n904_), .C2(G871), .ZN(G747));
  INV_X1    g0679(.A(G834), .ZN(new_n1109_));
  NAND2_X1  g0680(.A1(new_n1109_), .A2(new_n1106_), .ZN(new_n1110_));
  NOR2_X1   g0681(.A1(new_n902_), .A2(G20), .ZN(new_n1111_));
  OAI21_X1  g0682(.A(G4087), .B1(G76), .B2(G4088), .ZN(new_n1112_));
  OAI221_X1 g0683(.A(new_n1110_), .B1(new_n1111_), .B2(new_n1112_), .C1(G873), .C2(new_n904_), .ZN(G752));
  INV_X1    g0684(.A(G17), .ZN(new_n1114_));
  NAND2_X1  g0685(.A1(new_n1114_), .A2(G4088), .ZN(new_n1115_));
  OAI211_X1 g0686(.A(new_n1115_), .B(G4087), .C1(G73), .C2(G4088), .ZN(new_n1116_));
  OAI221_X1 g0687(.A(new_n1116_), .B1(new_n904_), .B2(G875), .C1(G836), .C2(new_n1107_), .ZN(G757));
  NAND2_X1  g0688(.A1(new_n872_), .A2(new_n898_), .ZN(new_n1118_));
  NOR2_X1   g0689(.A1(new_n902_), .A2(G70), .ZN(new_n1119_));
  OAI21_X1  g0690(.A(G4087), .B1(G67), .B2(G4088), .ZN(new_n1120_));
  OAI221_X1 g0691(.A(new_n1118_), .B1(new_n1119_), .B2(new_n1120_), .C1(G877), .C2(new_n904_), .ZN(G762));
  NOR2_X1   g0692(.A1(new_n938_), .A2(G4089), .ZN(new_n1122_));
  NAND2_X1  g0693(.A1(new_n918_), .A2(new_n1122_), .ZN(new_n1123_));
  XNOR2_X1  g0694(.A(new_n1123_), .B(KEYINPUT68), .ZN(new_n1124_));
  NOR2_X1   g0695(.A1(new_n939_), .A2(G37), .ZN(new_n1125_));
  OAI21_X1  g0696(.A(G4090), .B1(G43), .B2(G4089), .ZN(new_n1126_));
  OAI221_X1 g0697(.A(new_n1124_), .B1(new_n941_), .B2(G871), .C1(new_n1125_), .C2(new_n1126_), .ZN(G787));
  NAND2_X1  g0698(.A1(new_n1109_), .A2(new_n1122_), .ZN(new_n1128_));
  NOR2_X1   g0699(.A1(new_n939_), .A2(G20), .ZN(new_n1129_));
  OAI21_X1  g0700(.A(G4090), .B1(G76), .B2(G4089), .ZN(new_n1130_));
  OAI221_X1 g0701(.A(new_n1128_), .B1(new_n1129_), .B2(new_n1130_), .C1(G873), .C2(new_n941_), .ZN(G792));
  NAND2_X1  g0702(.A1(new_n1114_), .A2(G4089), .ZN(new_n1132_));
  OAI211_X1 g0703(.A(new_n1132_), .B(G4090), .C1(G73), .C2(G4089), .ZN(new_n1133_));
  INV_X1    g0704(.A(new_n1122_), .ZN(new_n1134_));
  OAI221_X1 g0705(.A(new_n1133_), .B1(new_n941_), .B2(G875), .C1(G836), .C2(new_n1134_), .ZN(G797));
  NAND2_X1  g0706(.A1(new_n872_), .A2(new_n936_), .ZN(new_n1136_));
  NOR2_X1   g0707(.A1(new_n939_), .A2(G70), .ZN(new_n1137_));
  OAI21_X1  g0708(.A(G4090), .B1(G67), .B2(G4089), .ZN(new_n1138_));
  OAI221_X1 g0709(.A(new_n1136_), .B1(new_n1137_), .B2(new_n1138_), .C1(G877), .C2(new_n941_), .ZN(new_n1139_));
  XNOR2_X1  g0710(.A(new_n1139_), .B(KEYINPUT69), .ZN(G802));
  INV_X1    g0711(.A(G871), .ZN(new_n1141_));
  NAND2_X1  g0712(.A1(new_n1141_), .A2(new_n1082_), .ZN(new_n1142_));
  NAND3_X1  g0713(.A1(G170), .A2(G1689), .A3(G1690), .ZN(new_n1143_));
  INV_X1    g0714(.A(G200), .ZN(new_n1144_));
  INV_X1    g0715(.A(G1690), .ZN(new_n1145_));
  OAI21_X1  g0716(.A(KEYINPUT70), .B1(new_n1144_), .B2(new_n1145_), .ZN(new_n1146_));
  NAND2_X1  g0717(.A1(new_n1146_), .A2(new_n1081_), .ZN(new_n1147_));
  NOR3_X1   g0718(.A1(new_n1144_), .A2(new_n1145_), .A3(KEYINPUT70), .ZN(new_n1148_));
  OAI21_X1  g0719(.A(new_n1143_), .B1(new_n1147_), .B2(new_n1148_), .ZN(new_n1149_));
  AOI21_X1  g0720(.A(new_n1149_), .B1(new_n918_), .B2(new_n1089_), .ZN(new_n1150_));
  AOI21_X1  g0721(.A(new_n1080_), .B1(new_n1142_), .B2(new_n1150_), .ZN(G642));
  OAI21_X1  g0722(.A(new_n1082_), .B1(new_n1000_), .B2(new_n1004_), .ZN(new_n1152_));
  OAI21_X1  g0723(.A(G1690), .B1(G188), .B2(G1689), .ZN(new_n1153_));
  INV_X1    g0724(.A(G158), .ZN(new_n1154_));
  AOI21_X1  g0725(.A(new_n1153_), .B1(new_n1154_), .B2(G1689), .ZN(new_n1155_));
  AOI21_X1  g0726(.A(new_n1155_), .B1(new_n872_), .B2(new_n1089_), .ZN(new_n1156_));
  AOI21_X1  g0727(.A(new_n1080_), .B1(new_n1152_), .B2(new_n1156_), .ZN(G664));
  INV_X1    g0728(.A(G836), .ZN(new_n1158_));
  NAND2_X1  g0729(.A1(new_n1158_), .A2(new_n1089_), .ZN(new_n1159_));
  OAI21_X1  g0730(.A(G1690), .B1(G155), .B2(G1689), .ZN(new_n1160_));
  INV_X1    g0731(.A(G152), .ZN(new_n1161_));
  AOI21_X1  g0732(.A(new_n1160_), .B1(new_n1161_), .B2(G1689), .ZN(new_n1162_));
  INV_X1    g0733(.A(G875), .ZN(new_n1163_));
  AOI21_X1  g0734(.A(new_n1162_), .B1(new_n1163_), .B2(new_n1082_), .ZN(new_n1164_));
  AOI21_X1  g0735(.A(new_n1080_), .B1(new_n1159_), .B2(new_n1164_), .ZN(G667));
  NAND2_X1  g0736(.A1(new_n982_), .A2(new_n1082_), .ZN(new_n1166_));
  XOR2_X1   g0737(.A(new_n1166_), .B(KEYINPUT71), .Z(new_n1167_));
  OAI21_X1  g0738(.A(G1690), .B1(G149), .B2(G1689), .ZN(new_n1168_));
  INV_X1    g0739(.A(G146), .ZN(new_n1169_));
  AOI21_X1  g0740(.A(new_n1168_), .B1(new_n1169_), .B2(G1689), .ZN(new_n1170_));
  AOI21_X1  g0741(.A(new_n1170_), .B1(new_n1109_), .B2(new_n1089_), .ZN(new_n1171_));
  AOI21_X1  g0742(.A(new_n1080_), .B1(new_n1167_), .B2(new_n1171_), .ZN(G670));
  NAND2_X1  g0743(.A1(new_n1141_), .A2(new_n1100_), .ZN(new_n1173_));
  NOR2_X1   g0744(.A1(new_n1096_), .A2(G170), .ZN(new_n1174_));
  AOI211_X1 g0745(.A(new_n1092_), .B(new_n1174_), .C1(new_n1144_), .C2(new_n1096_), .ZN(new_n1175_));
  NOR2_X1   g0746(.A1(G1691), .A2(G1694), .ZN(new_n1176_));
  AOI21_X1  g0747(.A(new_n1175_), .B1(new_n918_), .B2(new_n1176_), .ZN(new_n1177_));
  AOI21_X1  g0748(.A(new_n1080_), .B1(new_n1173_), .B2(new_n1177_), .ZN(G676));
  INV_X1    g0749(.A(new_n1100_), .ZN(new_n1179_));
  NOR2_X1   g0750(.A1(G877), .A2(new_n1179_), .ZN(new_n1180_));
  XNOR2_X1  g0751(.A(new_n1180_), .B(KEYINPUT72), .ZN(new_n1181_));
  OAI21_X1  g0752(.A(G1694), .B1(G188), .B2(G1691), .ZN(new_n1182_));
  AOI21_X1  g0753(.A(new_n1182_), .B1(new_n1154_), .B2(G1691), .ZN(new_n1183_));
  AOI21_X1  g0754(.A(new_n1183_), .B1(new_n872_), .B2(new_n1176_), .ZN(new_n1184_));
  AOI21_X1  g0755(.A(new_n1080_), .B1(new_n1181_), .B2(new_n1184_), .ZN(G696));
  NAND2_X1  g0756(.A1(new_n1158_), .A2(new_n1176_), .ZN(new_n1186_));
  OAI21_X1  g0757(.A(G1694), .B1(G155), .B2(G1691), .ZN(new_n1187_));
  AOI21_X1  g0758(.A(new_n1187_), .B1(new_n1161_), .B2(G1691), .ZN(new_n1188_));
  AOI21_X1  g0759(.A(new_n1188_), .B1(new_n1163_), .B2(new_n1100_), .ZN(new_n1189_));
  AOI21_X1  g0760(.A(new_n1080_), .B1(new_n1186_), .B2(new_n1189_), .ZN(G699));
  OAI21_X1  g0761(.A(G1694), .B1(G149), .B2(G1691), .ZN(new_n1191_));
  AOI21_X1  g0762(.A(new_n1191_), .B1(new_n1169_), .B2(G1691), .ZN(new_n1192_));
  AOI21_X1  g0763(.A(new_n1192_), .B1(new_n1109_), .B2(new_n1176_), .ZN(new_n1193_));
  NAND2_X1  g0764(.A1(new_n982_), .A2(new_n1100_), .ZN(new_n1194_));
  AOI21_X1  g0765(.A(new_n1080_), .B1(new_n1193_), .B2(new_n1194_), .ZN(G702));
  NAND2_X1  g0766(.A1(G135), .A2(G4115), .ZN(new_n1196_));
  NOR2_X1   g0767(.A1(new_n539_), .A2(G3717), .ZN(new_n1197_));
  INV_X1    g0768(.A(G3724), .ZN(new_n1198_));
  INV_X1    g0769(.A(G123), .ZN(new_n1199_));
  INV_X1    g0770(.A(G3717), .ZN(new_n1200_));
  OAI21_X1  g0771(.A(new_n1198_), .B1(new_n1199_), .B2(new_n1200_), .ZN(new_n1201_));
  OAI21_X1  g0772(.A(new_n1196_), .B1(new_n1197_), .B2(new_n1201_), .ZN(new_n1202_));
  NAND2_X1  g0773(.A1(new_n893_), .A2(G3717), .ZN(new_n1203_));
  XNOR2_X1  g0774(.A(new_n778_), .B(G132), .ZN(new_n1204_));
  AOI21_X1  g0775(.A(new_n1198_), .B1(new_n1204_), .B2(new_n1200_), .ZN(new_n1205_));
  AOI21_X1  g0776(.A(new_n1202_), .B1(new_n1203_), .B2(new_n1205_), .ZN(G818));
  XOR2_X1   g0777(.A(new_n893_), .B(new_n1204_), .Z(G813));
  NAND2_X1  g0778(.A1(new_n893_), .A2(new_n862_), .ZN(new_n1208_));
  AOI21_X1  g0779(.A(G4091), .B1(new_n1199_), .B2(G4092), .ZN(new_n1209_));
  OAI21_X1  g0780(.A(new_n1209_), .B1(new_n538_), .B2(G4092), .ZN(new_n1210_));
  NAND2_X1  g0781(.A1(new_n1208_), .A2(new_n1210_), .ZN(new_n1211_));
  INV_X1    g0782(.A(new_n1211_), .ZN(G824));
  AND2_X1   g0783(.A1(new_n1074_), .A2(new_n862_), .ZN(new_n1213_));
  OAI21_X1  g0784(.A(new_n861_), .B1(new_n854_), .B2(G121), .ZN(new_n1214_));
  AOI21_X1  g0785(.A(new_n1214_), .B1(new_n545_), .B2(new_n854_), .ZN(new_n1215_));
  NOR2_X1   g0786(.A1(new_n1213_), .A2(new_n1215_), .ZN(G826));
  NAND2_X1  g0787(.A1(new_n1068_), .A2(new_n862_), .ZN(new_n1217_));
  NAND2_X1  g0788(.A1(new_n534_), .A2(new_n854_), .ZN(new_n1218_));
  OAI211_X1 g0789(.A(new_n1218_), .B(new_n861_), .C1(G116), .C2(new_n854_), .ZN(new_n1219_));
  NAND2_X1  g0790(.A1(new_n1217_), .A2(new_n1219_), .ZN(new_n1220_));
  INV_X1    g0791(.A(new_n1220_), .ZN(G828));
  OAI21_X1  g0792(.A(new_n861_), .B1(new_n854_), .B2(G112), .ZN(new_n1222_));
  AOI21_X1  g0793(.A(new_n1222_), .B1(new_n528_), .B2(new_n854_), .ZN(new_n1223_));
  AOI21_X1  g0794(.A(new_n1223_), .B1(new_n1071_), .B2(new_n862_), .ZN(new_n1224_));
  XNOR2_X1  g0795(.A(new_n1224_), .B(KEYINPUT73), .ZN(new_n1225_));
  INV_X1    g0796(.A(new_n1225_), .ZN(G830));
  NAND3_X1  g0797(.A1(G601), .A2(G245), .A3(G559), .ZN(new_n1227_));
  OR3_X1    g0798(.A1(G1002), .A2(G847), .A3(new_n1227_), .ZN(new_n1228_));
  NOR4_X1   g0799(.A1(G1000), .A2(G998), .A3(G1004), .A4(new_n1228_), .ZN(G854));
  OR2_X1    g0800(.A1(new_n1047_), .A2(new_n863_), .ZN(new_n1230_));
  NAND2_X1  g0801(.A1(new_n593_), .A2(new_n854_), .ZN(new_n1231_));
  OAI211_X1 g0802(.A(new_n1231_), .B(new_n861_), .C1(G115), .C2(new_n854_), .ZN(new_n1232_));
  NAND2_X1  g0803(.A1(new_n1230_), .A2(new_n1232_), .ZN(new_n1233_));
  INV_X1    g0804(.A(new_n1233_), .ZN(G863));
  AOI21_X1  g0805(.A(new_n863_), .B1(new_n1052_), .B2(new_n1054_), .ZN(new_n1235_));
  OAI21_X1  g0806(.A(new_n861_), .B1(new_n854_), .B2(G114), .ZN(new_n1236_));
  AOI21_X1  g0807(.A(new_n1236_), .B1(new_n628_), .B2(new_n854_), .ZN(new_n1237_));
  NOR2_X1   g0808(.A1(new_n1235_), .A2(new_n1237_), .ZN(G865));
  NAND2_X1  g0809(.A1(new_n1058_), .A2(new_n862_), .ZN(new_n1239_));
  OR2_X1    g0810(.A1(new_n1239_), .A2(KEYINPUT74), .ZN(new_n1240_));
  NAND2_X1  g0811(.A1(new_n610_), .A2(new_n854_), .ZN(new_n1241_));
  OAI211_X1 g0812(.A(new_n1241_), .B(new_n861_), .C1(G53), .C2(new_n854_), .ZN(new_n1242_));
  NAND2_X1  g0813(.A1(new_n1239_), .A2(KEYINPUT74), .ZN(new_n1243_));
  NAND3_X1  g0814(.A1(new_n1240_), .A2(new_n1242_), .A3(new_n1243_), .ZN(new_n1244_));
  INV_X1    g0815(.A(new_n1244_), .ZN(G867));
  NAND2_X1  g0816(.A1(new_n616_), .A2(new_n854_), .ZN(new_n1246_));
  OAI211_X1 g0817(.A(new_n1246_), .B(new_n861_), .C1(G113), .C2(new_n854_), .ZN(new_n1247_));
  OAI21_X1  g0818(.A(new_n1247_), .B1(new_n1049_), .B2(new_n863_), .ZN(new_n1248_));
  XNOR2_X1  g0819(.A(new_n1248_), .B(KEYINPUT75), .ZN(new_n1249_));
  INV_X1    g0820(.A(new_n1249_), .ZN(G869));
  NAND3_X1  g0821(.A1(new_n939_), .A2(G109), .A3(G4090), .ZN(new_n1251_));
  XNOR2_X1  g0822(.A(new_n1251_), .B(KEYINPUT76), .ZN(new_n1252_));
  AND3_X1   g0823(.A1(G106), .A2(G4089), .A3(G4090), .ZN(new_n1253_));
  AOI211_X1 g0824(.A(new_n1252_), .B(new_n1253_), .C1(new_n1233_), .C2(new_n940_), .ZN(new_n1254_));
  OAI21_X1  g0825(.A(new_n1254_), .B1(G824), .B2(new_n1134_), .ZN(G712));
  OR2_X1    g0826(.A1(G109), .A2(G4088), .ZN(new_n1256_));
  OAI211_X1 g0827(.A(new_n1256_), .B(G4087), .C1(G106), .C2(new_n902_), .ZN(new_n1257_));
  OAI221_X1 g0828(.A(new_n1257_), .B1(new_n904_), .B2(G863), .C1(G824), .C2(new_n1107_), .ZN(G727));
  OAI21_X1  g0829(.A(G4087), .B1(G46), .B2(G4088), .ZN(new_n1259_));
  INV_X1    g0830(.A(G49), .ZN(new_n1260_));
  AOI21_X1  g0831(.A(new_n1259_), .B1(new_n1260_), .B2(G4088), .ZN(new_n1261_));
  INV_X1    g0832(.A(G865), .ZN(new_n1262_));
  AOI21_X1  g0833(.A(new_n1261_), .B1(new_n1262_), .B2(new_n903_), .ZN(new_n1263_));
  OAI21_X1  g0834(.A(new_n1263_), .B1(G826), .B2(new_n1107_), .ZN(G732));
  INV_X1    g0835(.A(G103), .ZN(new_n1265_));
  NAND2_X1  g0836(.A1(new_n1265_), .A2(G4088), .ZN(new_n1266_));
  OAI211_X1 g0837(.A(new_n1266_), .B(G4087), .C1(G100), .C2(G4088), .ZN(new_n1267_));
  OAI221_X1 g0838(.A(new_n1267_), .B1(new_n1107_), .B2(G828), .C1(G867), .C2(new_n904_), .ZN(G737));
  OAI21_X1  g0839(.A(G4087), .B1(G91), .B2(G4088), .ZN(new_n1269_));
  INV_X1    g0840(.A(G40), .ZN(new_n1270_));
  AOI21_X1  g0841(.A(new_n1269_), .B1(new_n1270_), .B2(G4088), .ZN(new_n1271_));
  AOI21_X1  g0842(.A(new_n1271_), .B1(new_n1249_), .B2(new_n903_), .ZN(new_n1272_));
  OAI21_X1  g0843(.A(new_n1272_), .B1(G830), .B2(new_n1107_), .ZN(G742));
  OAI21_X1  g0844(.A(G4090), .B1(G46), .B2(G4089), .ZN(new_n1274_));
  AOI21_X1  g0845(.A(new_n1274_), .B1(new_n1260_), .B2(G4089), .ZN(new_n1275_));
  AOI21_X1  g0846(.A(new_n1275_), .B1(new_n1262_), .B2(new_n940_), .ZN(new_n1276_));
  OAI21_X1  g0847(.A(new_n1276_), .B1(G826), .B2(new_n1134_), .ZN(G772));
  NAND2_X1  g0848(.A1(new_n1265_), .A2(G4089), .ZN(new_n1278_));
  OAI211_X1 g0849(.A(new_n1278_), .B(G4090), .C1(G100), .C2(G4089), .ZN(new_n1279_));
  OAI221_X1 g0850(.A(new_n1279_), .B1(new_n1134_), .B2(G828), .C1(G867), .C2(new_n941_), .ZN(G777));
  OAI21_X1  g0851(.A(G4090), .B1(G91), .B2(G4089), .ZN(new_n1281_));
  AOI21_X1  g0852(.A(new_n1281_), .B1(new_n1270_), .B2(G4089), .ZN(new_n1282_));
  AOI21_X1  g0853(.A(new_n1282_), .B1(new_n1249_), .B2(new_n940_), .ZN(new_n1283_));
  OAI21_X1  g0854(.A(new_n1283_), .B1(G830), .B2(new_n1134_), .ZN(G782));
  NAND2_X1  g0855(.A1(new_n1225_), .A2(new_n1089_), .ZN(new_n1285_));
  OAI21_X1  g0856(.A(G1690), .B1(G203), .B2(G1689), .ZN(new_n1286_));
  INV_X1    g0857(.A(G173), .ZN(new_n1287_));
  AOI21_X1  g0858(.A(new_n1286_), .B1(new_n1287_), .B2(G1689), .ZN(new_n1288_));
  AOI21_X1  g0859(.A(new_n1288_), .B1(new_n1249_), .B2(new_n1082_), .ZN(new_n1289_));
  AOI21_X1  g0860(.A(new_n1080_), .B1(new_n1285_), .B2(new_n1289_), .ZN(G645));
  OAI21_X1  g0861(.A(G1690), .B1(G197), .B2(G1689), .ZN(new_n1291_));
  INV_X1    g0862(.A(G167), .ZN(new_n1292_));
  AOI21_X1  g0863(.A(new_n1291_), .B1(new_n1292_), .B2(G1689), .ZN(new_n1293_));
  AOI21_X1  g0864(.A(new_n1293_), .B1(new_n1244_), .B2(new_n1082_), .ZN(new_n1294_));
  NAND2_X1  g0865(.A1(new_n1220_), .A2(new_n1089_), .ZN(new_n1295_));
  AOI21_X1  g0866(.A(new_n1080_), .B1(new_n1294_), .B2(new_n1295_), .ZN(G648));
  OAI21_X1  g0867(.A(new_n1089_), .B1(new_n1213_), .B2(new_n1215_), .ZN(new_n1297_));
  OAI21_X1  g0868(.A(G1690), .B1(G194), .B2(G1689), .ZN(new_n1298_));
  INV_X1    g0869(.A(G164), .ZN(new_n1299_));
  AOI21_X1  g0870(.A(new_n1298_), .B1(new_n1299_), .B2(G1689), .ZN(new_n1300_));
  AOI21_X1  g0871(.A(new_n1300_), .B1(new_n1262_), .B2(new_n1082_), .ZN(new_n1301_));
  AOI21_X1  g0872(.A(new_n1080_), .B1(new_n1297_), .B2(new_n1301_), .ZN(G651));
  NAND2_X1  g0873(.A1(new_n1211_), .A2(new_n1089_), .ZN(new_n1303_));
  OAI21_X1  g0874(.A(G1690), .B1(G191), .B2(G1689), .ZN(new_n1304_));
  INV_X1    g0875(.A(G161), .ZN(new_n1305_));
  AOI21_X1  g0876(.A(new_n1304_), .B1(new_n1305_), .B2(G1689), .ZN(new_n1306_));
  AOI21_X1  g0877(.A(new_n1306_), .B1(new_n1233_), .B2(new_n1082_), .ZN(new_n1307_));
  AOI21_X1  g0878(.A(new_n1080_), .B1(new_n1303_), .B2(new_n1307_), .ZN(G654));
  NAND2_X1  g0879(.A1(new_n1225_), .A2(new_n1176_), .ZN(new_n1309_));
  OAI21_X1  g0880(.A(G1694), .B1(G203), .B2(G1691), .ZN(new_n1310_));
  AOI21_X1  g0881(.A(new_n1310_), .B1(new_n1287_), .B2(G1691), .ZN(new_n1311_));
  XNOR2_X1  g0882(.A(new_n1311_), .B(KEYINPUT77), .ZN(new_n1312_));
  AOI21_X1  g0883(.A(new_n1312_), .B1(new_n1249_), .B2(new_n1100_), .ZN(new_n1313_));
  AOI21_X1  g0884(.A(new_n1080_), .B1(new_n1309_), .B2(new_n1313_), .ZN(G679));
  NAND2_X1  g0885(.A1(new_n1220_), .A2(new_n1176_), .ZN(new_n1315_));
  NAND2_X1  g0886(.A1(new_n1292_), .A2(G1691), .ZN(new_n1316_));
  OAI211_X1 g0887(.A(new_n1316_), .B(G1694), .C1(G197), .C2(G1691), .ZN(new_n1317_));
  OAI211_X1 g0888(.A(new_n1315_), .B(new_n1317_), .C1(G867), .C2(new_n1179_), .ZN(new_n1318_));
  NAND2_X1  g0889(.A1(new_n1318_), .A2(G137), .ZN(new_n1319_));
  XNOR2_X1  g0890(.A(new_n1319_), .B(KEYINPUT78), .ZN(G682));
  OAI21_X1  g0891(.A(new_n1176_), .B1(new_n1213_), .B2(new_n1215_), .ZN(new_n1321_));
  NAND2_X1  g0892(.A1(new_n1299_), .A2(G1691), .ZN(new_n1322_));
  OAI211_X1 g0893(.A(new_n1322_), .B(G1694), .C1(G194), .C2(G1691), .ZN(new_n1323_));
  NAND3_X1  g0894(.A1(new_n1321_), .A2(KEYINPUT79), .A3(new_n1323_), .ZN(new_n1324_));
  OAI21_X1  g0895(.A(new_n1324_), .B1(new_n1179_), .B2(G865), .ZN(new_n1325_));
  AOI21_X1  g0896(.A(KEYINPUT79), .B1(new_n1321_), .B2(new_n1323_), .ZN(new_n1326_));
  OAI21_X1  g0897(.A(G137), .B1(new_n1325_), .B2(new_n1326_), .ZN(new_n1327_));
  XNOR2_X1  g0898(.A(new_n1327_), .B(KEYINPUT80), .ZN(G685));
  NOR2_X1   g0899(.A1(G824), .A2(G1694), .ZN(new_n1329_));
  AOI21_X1  g0900(.A(G1691), .B1(new_n1329_), .B2(KEYINPUT81), .ZN(new_n1330_));
  OAI21_X1  g0901(.A(new_n1330_), .B1(KEYINPUT81), .B2(new_n1329_), .ZN(new_n1331_));
  NAND2_X1  g0902(.A1(new_n1305_), .A2(G1691), .ZN(new_n1332_));
  OAI211_X1 g0903(.A(new_n1332_), .B(G1694), .C1(G191), .C2(G1691), .ZN(new_n1333_));
  NOR2_X1   g0904(.A1(G863), .A2(new_n1179_), .ZN(new_n1334_));
  OAI21_X1  g0905(.A(new_n1333_), .B1(new_n1334_), .B2(KEYINPUT82), .ZN(new_n1335_));
  AOI21_X1  g0906(.A(new_n1335_), .B1(KEYINPUT82), .B2(new_n1334_), .ZN(new_n1336_));
  AOI21_X1  g0907(.A(new_n1080_), .B1(new_n1331_), .B2(new_n1336_), .ZN(G688));
  OAI21_X1  g0908(.A(G4092), .B1(G120), .B2(G4091), .ZN(new_n1338_));
  XOR2_X1   g0909(.A(new_n1338_), .B(KEYINPUT98), .Z(new_n1339_));
  NAND3_X1  g0910(.A1(G248), .A2(G324), .A3(G503), .ZN(new_n1340_));
  XNOR2_X1  g0911(.A(new_n1340_), .B(KEYINPUT95), .ZN(new_n1341_));
  NAND2_X1  g0912(.A1(new_n503_), .A2(G251), .ZN(new_n1342_));
  AOI21_X1  g0913(.A(G503), .B1(new_n499_), .B2(G254), .ZN(new_n1343_));
  OAI21_X1  g0914(.A(new_n1343_), .B1(new_n524_), .B2(new_n499_), .ZN(new_n1344_));
  NAND3_X1  g0915(.A1(new_n1341_), .A2(new_n1342_), .A3(new_n1344_), .ZN(new_n1345_));
  XNOR2_X1  g0916(.A(new_n1345_), .B(KEYINPUT96), .ZN(new_n1346_));
  MUX2_X1   g0917(.A(new_n524_), .B(G248), .S(G514), .Z(new_n1347_));
  XNOR2_X1  g0918(.A(new_n1346_), .B(new_n1347_), .ZN(new_n1348_));
  OR2_X1    g0919(.A1(new_n1348_), .A2(new_n547_), .ZN(new_n1349_));
  NAND3_X1  g0920(.A1(new_n508_), .A2(G251), .A3(G523), .ZN(new_n1350_));
  XNOR2_X1  g0921(.A(new_n1350_), .B(KEYINPUT93), .ZN(new_n1351_));
  NAND3_X1  g0922(.A1(G248), .A2(G341), .A3(G523), .ZN(new_n1352_));
  NOR2_X1   g0923(.A1(new_n524_), .A2(new_n508_), .ZN(new_n1353_));
  OAI21_X1  g0924(.A(new_n732_), .B1(new_n537_), .B2(G341), .ZN(new_n1354_));
  OAI211_X1 g0925(.A(new_n1351_), .B(new_n1352_), .C1(new_n1353_), .C2(new_n1354_), .ZN(new_n1355_));
  XOR2_X1   g0926(.A(new_n1355_), .B(KEYINPUT94), .Z(new_n1356_));
  OAI21_X1  g0927(.A(new_n743_), .B1(new_n537_), .B2(G351), .ZN(new_n1357_));
  AOI21_X1  g0928(.A(new_n1357_), .B1(G242), .B2(G351), .ZN(new_n1358_));
  INV_X1    g0929(.A(G248), .ZN(new_n1359_));
  OAI22_X1  g0930(.A1(new_n515_), .A2(new_n544_), .B1(new_n1359_), .B2(new_n516_), .ZN(new_n1360_));
  AOI21_X1  g0931(.A(new_n1358_), .B1(new_n1360_), .B2(G534), .ZN(new_n1361_));
  XNOR2_X1  g0932(.A(new_n1356_), .B(new_n1361_), .ZN(new_n1362_));
  NOR2_X1   g0933(.A1(new_n1349_), .A2(new_n1362_), .ZN(new_n1363_));
  XNOR2_X1  g0934(.A(new_n1363_), .B(KEYINPUT97), .ZN(new_n1364_));
  NAND2_X1  g0935(.A1(new_n1348_), .A2(new_n547_), .ZN(new_n1365_));
  NAND3_X1  g0936(.A1(new_n1349_), .A2(new_n1362_), .A3(new_n1365_), .ZN(new_n1366_));
  OAI211_X1 g0937(.A(new_n1364_), .B(new_n1366_), .C1(new_n1362_), .C2(new_n1365_), .ZN(new_n1367_));
  XNOR2_X1  g0938(.A(new_n528_), .B(new_n534_), .ZN(new_n1368_));
  XNOR2_X1  g0939(.A(new_n545_), .B(new_n538_), .ZN(new_n1369_));
  XNOR2_X1  g0940(.A(new_n1368_), .B(new_n1369_), .ZN(new_n1370_));
  XNOR2_X1  g0941(.A(new_n1367_), .B(new_n1370_), .ZN(new_n1371_));
  AOI21_X1  g0942(.A(new_n1339_), .B1(new_n1371_), .B2(new_n857_), .ZN(new_n1372_));
  NAND3_X1  g0943(.A1(new_n738_), .A2(G2174), .A3(new_n756_), .ZN(new_n1373_));
  NAND2_X1  g0944(.A1(new_n765_), .A2(new_n1069_), .ZN(new_n1374_));
  NAND2_X1  g0945(.A1(new_n771_), .A2(new_n1374_), .ZN(new_n1375_));
  XNOR2_X1  g0946(.A(new_n839_), .B(new_n1375_), .ZN(new_n1376_));
  OAI21_X1  g0947(.A(new_n837_), .B1(new_n766_), .B2(new_n836_), .ZN(new_n1377_));
  NOR2_X1   g0948(.A1(new_n761_), .A2(new_n764_), .ZN(new_n1378_));
  OAI211_X1 g0949(.A(new_n1377_), .B(KEYINPUT90), .C1(new_n1378_), .C2(new_n837_), .ZN(new_n1379_));
  OAI21_X1  g0950(.A(new_n1379_), .B1(KEYINPUT90), .B2(new_n1377_), .ZN(new_n1380_));
  XNOR2_X1  g0951(.A(new_n1376_), .B(new_n1380_), .ZN(new_n1381_));
  INV_X1    g0952(.A(new_n778_), .ZN(new_n1382_));
  NOR2_X1   g0953(.A1(new_n1381_), .A2(new_n1382_), .ZN(new_n1383_));
  XNOR2_X1  g0954(.A(new_n1383_), .B(KEYINPUT91), .ZN(new_n1384_));
  NAND2_X1  g0955(.A1(new_n1381_), .A2(new_n779_), .ZN(new_n1385_));
  XOR2_X1   g0956(.A(new_n1385_), .B(KEYINPUT92), .Z(new_n1386_));
  OAI211_X1 g0957(.A(new_n850_), .B(new_n1373_), .C1(new_n1384_), .C2(new_n1386_), .ZN(new_n1387_));
  NAND2_X1  g0958(.A1(new_n850_), .A2(new_n1373_), .ZN(new_n1388_));
  XNOR2_X1  g0959(.A(new_n887_), .B(new_n1069_), .ZN(new_n1389_));
  NAND2_X1  g0960(.A1(new_n886_), .A2(new_n763_), .ZN(new_n1390_));
  OAI21_X1  g0961(.A(new_n1390_), .B1(new_n1378_), .B2(new_n886_), .ZN(new_n1391_));
  XNOR2_X1  g0962(.A(new_n1389_), .B(new_n1391_), .ZN(new_n1392_));
  NAND2_X1  g0963(.A1(new_n1392_), .A2(new_n1382_), .ZN(new_n1393_));
  OAI211_X1 g0964(.A(new_n1388_), .B(new_n1393_), .C1(new_n779_), .C2(new_n1392_), .ZN(new_n1394_));
  NAND2_X1  g0965(.A1(new_n1387_), .A2(new_n1394_), .ZN(new_n1395_));
  NAND2_X1  g0966(.A1(new_n1395_), .A2(new_n1073_), .ZN(new_n1396_));
  NAND3_X1  g0967(.A1(new_n1387_), .A2(new_n775_), .A3(new_n1394_), .ZN(new_n1397_));
  NAND2_X1  g0968(.A1(new_n1396_), .A2(new_n1397_), .ZN(new_n1398_));
  NOR2_X1   g0969(.A1(new_n910_), .A2(KEYINPUT88), .ZN(new_n1399_));
  MUX2_X1   g0970(.A(new_n1399_), .B(new_n733_), .S(new_n842_), .Z(new_n1400_));
  NAND3_X1  g0971(.A1(new_n751_), .A2(new_n736_), .A3(new_n728_), .ZN(new_n1401_));
  AND2_X1   g0972(.A1(new_n1401_), .A2(new_n911_), .ZN(new_n1402_));
  XNOR2_X1  g0973(.A(new_n1400_), .B(new_n1402_), .ZN(new_n1403_));
  XNOR2_X1  g0974(.A(new_n751_), .B(new_n755_), .ZN(new_n1404_));
  XNOR2_X1  g0975(.A(new_n1403_), .B(new_n1404_), .ZN(new_n1405_));
  OR2_X1    g0976(.A1(new_n1405_), .A2(new_n720_), .ZN(new_n1406_));
  NAND2_X1  g0977(.A1(new_n1405_), .A2(new_n720_), .ZN(new_n1407_));
  AOI21_X1  g0978(.A(new_n727_), .B1(new_n1406_), .B2(new_n1407_), .ZN(new_n1408_));
  INV_X1    g0979(.A(new_n1408_), .ZN(new_n1409_));
  INV_X1    g0980(.A(KEYINPUT89), .ZN(new_n1410_));
  NAND2_X1  g0981(.A1(new_n1407_), .A2(new_n1410_), .ZN(new_n1411_));
  NAND3_X1  g0982(.A1(new_n1406_), .A2(new_n727_), .A3(new_n1407_), .ZN(new_n1412_));
  NAND4_X1  g0983(.A1(new_n1409_), .A2(new_n736_), .A3(new_n1411_), .A4(new_n1412_), .ZN(new_n1413_));
  NAND2_X1  g0984(.A1(new_n1411_), .A2(new_n736_), .ZN(new_n1414_));
  INV_X1    g0985(.A(new_n1412_), .ZN(new_n1415_));
  OAI21_X1  g0986(.A(new_n1414_), .B1(new_n1415_), .B2(new_n1408_), .ZN(new_n1416_));
  NAND3_X1  g0987(.A1(new_n1413_), .A2(new_n1416_), .A3(G2174), .ZN(new_n1417_));
  INV_X1    g0988(.A(new_n1417_), .ZN(new_n1418_));
  AND2_X1   g0989(.A1(new_n842_), .A2(new_n844_), .ZN(new_n1419_));
  AOI21_X1  g0990(.A(new_n843_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n1420_));
  NAND3_X1  g0991(.A1(new_n909_), .A2(new_n846_), .A3(new_n843_), .ZN(new_n1421_));
  INV_X1    g0992(.A(new_n1421_), .ZN(new_n1422_));
  OAI21_X1  g0993(.A(new_n1419_), .B1(new_n1420_), .B2(new_n1422_), .ZN(new_n1423_));
  INV_X1    g0994(.A(KEYINPUT83), .ZN(new_n1424_));
  NAND2_X1  g0995(.A1(new_n1421_), .A2(new_n1424_), .ZN(new_n1425_));
  NAND4_X1  g0996(.A1(new_n909_), .A2(new_n846_), .A3(KEYINPUT83), .A4(new_n843_), .ZN(new_n1426_));
  OAI211_X1 g0997(.A(new_n733_), .B(new_n755_), .C1(new_n735_), .C2(new_n925_), .ZN(new_n1427_));
  NAND3_X1  g0998(.A1(new_n1425_), .A2(new_n1426_), .A3(new_n1427_), .ZN(new_n1428_));
  AOI21_X1  g0999(.A(new_n1428_), .B1(new_n844_), .B2(new_n842_), .ZN(new_n1429_));
  INV_X1    g1000(.A(new_n1429_), .ZN(new_n1430_));
  AND3_X1   g1001(.A1(new_n1423_), .A2(new_n913_), .A3(new_n1430_), .ZN(new_n1431_));
  AND3_X1   g1002(.A1(new_n1428_), .A2(new_n844_), .A3(new_n842_), .ZN(new_n1432_));
  OAI21_X1  g1003(.A(new_n912_), .B1(new_n1432_), .B2(new_n1429_), .ZN(new_n1433_));
  INV_X1    g1004(.A(KEYINPUT84), .ZN(new_n1434_));
  NAND2_X1  g1005(.A1(new_n1433_), .A2(new_n1434_), .ZN(new_n1435_));
  OAI211_X1 g1006(.A(KEYINPUT84), .B(new_n912_), .C1(new_n1432_), .C2(new_n1429_), .ZN(new_n1436_));
  NAND2_X1  g1007(.A1(new_n1435_), .A2(new_n1436_), .ZN(new_n1437_));
  OAI21_X1  g1008(.A(new_n755_), .B1(new_n1431_), .B2(new_n1437_), .ZN(new_n1438_));
  NAND3_X1  g1009(.A1(new_n1423_), .A2(new_n913_), .A3(new_n1430_), .ZN(new_n1439_));
  NAND4_X1  g1010(.A1(new_n1439_), .A2(new_n843_), .A3(new_n1435_), .A4(new_n1436_), .ZN(new_n1440_));
  NAND3_X1  g1011(.A1(new_n1438_), .A2(KEYINPUT85), .A3(new_n1440_), .ZN(new_n1441_));
  INV_X1    g1012(.A(KEYINPUT85), .ZN(new_n1442_));
  OAI211_X1 g1013(.A(new_n1442_), .B(new_n755_), .C1(new_n1431_), .C2(new_n1437_), .ZN(new_n1443_));
  NAND3_X1  g1014(.A1(new_n1441_), .A2(new_n752_), .A3(new_n1443_), .ZN(new_n1444_));
  OR2_X1    g1015(.A1(new_n1432_), .A2(new_n1429_), .ZN(new_n1445_));
  AOI21_X1  g1016(.A(new_n843_), .B1(new_n1445_), .B2(new_n1402_), .ZN(new_n1446_));
  NAND2_X1  g1017(.A1(new_n1423_), .A2(new_n1430_), .ZN(new_n1447_));
  OAI21_X1  g1018(.A(new_n1446_), .B1(new_n1447_), .B2(new_n913_), .ZN(new_n1448_));
  NAND2_X1  g1019(.A1(new_n1448_), .A2(KEYINPUT86), .ZN(new_n1449_));
  INV_X1    g1020(.A(KEYINPUT86), .ZN(new_n1450_));
  OAI211_X1 g1021(.A(new_n1446_), .B(new_n1450_), .C1(new_n1447_), .C2(new_n913_), .ZN(new_n1451_));
  NAND4_X1  g1022(.A1(new_n1449_), .A2(new_n751_), .A3(new_n1440_), .A4(new_n1451_), .ZN(new_n1452_));
  NAND3_X1  g1023(.A1(new_n1444_), .A2(new_n719_), .A3(new_n1452_), .ZN(new_n1453_));
  NAND3_X1  g1024(.A1(new_n1441_), .A2(new_n751_), .A3(new_n1443_), .ZN(new_n1454_));
  NAND4_X1  g1025(.A1(new_n1449_), .A2(new_n752_), .A3(new_n1440_), .A4(new_n1451_), .ZN(new_n1455_));
  NAND3_X1  g1026(.A1(new_n1454_), .A2(new_n720_), .A3(new_n1455_), .ZN(new_n1456_));
  NAND3_X1  g1027(.A1(new_n1453_), .A2(new_n1456_), .A3(new_n736_), .ZN(new_n1457_));
  AND3_X1   g1028(.A1(new_n1444_), .A2(new_n719_), .A3(new_n1452_), .ZN(new_n1458_));
  AOI21_X1  g1029(.A(new_n719_), .B1(new_n1444_), .B2(new_n1452_), .ZN(new_n1459_));
  NOR2_X1   g1030(.A1(new_n1458_), .A2(new_n1459_), .ZN(new_n1460_));
  OAI211_X1 g1031(.A(new_n728_), .B(new_n1457_), .C1(new_n1460_), .C2(new_n736_), .ZN(new_n1461_));
  INV_X1    g1032(.A(G2174), .ZN(new_n1462_));
  AND2_X1   g1033(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1463_));
  NAND2_X1  g1034(.A1(new_n1453_), .A2(new_n1456_), .ZN(new_n1464_));
  INV_X1    g1035(.A(new_n736_), .ZN(new_n1465_));
  NAND2_X1  g1036(.A1(new_n1464_), .A2(new_n1465_), .ZN(new_n1466_));
  NAND2_X1  g1037(.A1(new_n1444_), .A2(new_n1452_), .ZN(new_n1467_));
  NAND2_X1  g1038(.A1(new_n1467_), .A2(new_n720_), .ZN(new_n1468_));
  NAND3_X1  g1039(.A1(new_n1468_), .A2(new_n736_), .A3(new_n1453_), .ZN(new_n1469_));
  NAND3_X1  g1040(.A1(new_n1466_), .A2(new_n1469_), .A3(KEYINPUT87), .ZN(new_n1470_));
  INV_X1    g1041(.A(KEYINPUT87), .ZN(new_n1471_));
  NAND4_X1  g1042(.A1(new_n1468_), .A2(new_n1471_), .A3(new_n736_), .A4(new_n1453_), .ZN(new_n1472_));
  NAND3_X1  g1043(.A1(new_n1470_), .A2(new_n727_), .A3(new_n1472_), .ZN(new_n1473_));
  AOI211_X1 g1044(.A(new_n1398_), .B(new_n1418_), .C1(new_n1463_), .C2(new_n1473_), .ZN(new_n1474_));
  INV_X1    g1045(.A(new_n1398_), .ZN(new_n1475_));
  AND3_X1   g1046(.A1(new_n1466_), .A2(new_n1469_), .A3(KEYINPUT87), .ZN(new_n1476_));
  NAND2_X1  g1047(.A1(new_n1472_), .A2(new_n727_), .ZN(new_n1477_));
  OAI211_X1 g1048(.A(new_n1462_), .B(new_n1461_), .C1(new_n1476_), .C2(new_n1477_), .ZN(new_n1478_));
  AOI21_X1  g1049(.A(new_n1475_), .B1(new_n1478_), .B2(new_n1417_), .ZN(new_n1479_));
  NOR2_X1   g1050(.A1(new_n1474_), .A2(new_n1479_), .ZN(new_n1480_));
  INV_X1    g1051(.A(new_n1480_), .ZN(new_n1481_));
  OAI21_X1  g1052(.A(new_n1372_), .B1(new_n1481_), .B2(new_n863_), .ZN(G843));
  OAI21_X1  g1053(.A(G4092), .B1(G118), .B2(G4091), .ZN(new_n1483_));
  NOR2_X1   g1054(.A1(new_n606_), .A2(new_n1359_), .ZN(new_n1484_));
  XNOR2_X1  g1055(.A(new_n1484_), .B(KEYINPUT119), .ZN(new_n1485_));
  AOI21_X1  g1056(.A(G468), .B1(G218), .B2(G242), .ZN(new_n1486_));
  INV_X1    g1057(.A(new_n1486_), .ZN(new_n1487_));
  OAI22_X1  g1058(.A1(new_n1487_), .A2(KEYINPUT118), .B1(G218), .B2(new_n537_), .ZN(new_n1488_));
  AND2_X1   g1059(.A1(new_n1487_), .A2(KEYINPUT118), .ZN(new_n1489_));
  OAI221_X1 g1060(.A(new_n1485_), .B1(new_n1488_), .B2(new_n1489_), .C1(new_n544_), .C2(new_n609_), .ZN(new_n1490_));
  XOR2_X1   g1061(.A(new_n592_), .B(new_n1490_), .Z(new_n1491_));
  NAND2_X1  g1062(.A1(G234), .A2(G242), .ZN(new_n1492_));
  OAI211_X1 g1063(.A(new_n1492_), .B(new_n594_), .C1(G234), .C2(new_n537_), .ZN(new_n1493_));
  OAI221_X1 g1064(.A(new_n1493_), .B1(new_n1359_), .B2(new_n597_), .C1(new_n595_), .C2(new_n544_), .ZN(new_n1494_));
  XNOR2_X1  g1065(.A(new_n1491_), .B(new_n1494_), .ZN(new_n1495_));
  OAI21_X1  g1066(.A(new_n619_), .B1(new_n623_), .B2(new_n524_), .ZN(new_n1496_));
  OR2_X1    g1067(.A1(new_n1496_), .A2(KEYINPUT120), .ZN(new_n1497_));
  NAND2_X1  g1068(.A1(new_n1496_), .A2(KEYINPUT120), .ZN(new_n1498_));
  OAI211_X1 g1069(.A(new_n1497_), .B(new_n1498_), .C1(G210), .C2(new_n537_), .ZN(new_n1499_));
  AOI22_X1  g1070(.A1(new_n621_), .A2(G251), .B1(G210), .B2(G248), .ZN(new_n1500_));
  OAI21_X1  g1071(.A(new_n1499_), .B1(new_n619_), .B2(new_n1500_), .ZN(new_n1501_));
  OAI21_X1  g1072(.A(new_n576_), .B1(new_n537_), .B2(G265), .ZN(new_n1502_));
  NOR2_X1   g1073(.A1(new_n524_), .A2(new_n577_), .ZN(new_n1503_));
  NOR2_X1   g1074(.A1(new_n577_), .A2(G248), .ZN(new_n1504_));
  OAI21_X1  g1075(.A(G400), .B1(G251), .B2(G265), .ZN(new_n1505_));
  OAI22_X1  g1076(.A1(new_n1502_), .A2(new_n1503_), .B1(new_n1504_), .B2(new_n1505_), .ZN(new_n1506_));
  XNOR2_X1  g1077(.A(new_n1501_), .B(new_n1506_), .ZN(new_n1507_));
  NAND3_X1  g1078(.A1(new_n562_), .A2(G251), .A3(G389), .ZN(new_n1508_));
  XOR2_X1   g1079(.A(new_n1508_), .B(KEYINPUT114), .Z(new_n1509_));
  NAND3_X1  g1080(.A1(G248), .A2(G257), .A3(G389), .ZN(new_n1510_));
  NOR2_X1   g1081(.A1(new_n524_), .A2(new_n562_), .ZN(new_n1511_));
  OAI21_X1  g1082(.A(new_n561_), .B1(new_n537_), .B2(G257), .ZN(new_n1512_));
  OAI211_X1 g1083(.A(new_n1509_), .B(new_n1510_), .C1(new_n1511_), .C2(new_n1512_), .ZN(new_n1513_));
  XOR2_X1   g1084(.A(new_n1507_), .B(new_n1513_), .Z(new_n1514_));
  XNOR2_X1  g1085(.A(new_n1495_), .B(new_n1514_), .ZN(new_n1515_));
  OAI21_X1  g1086(.A(new_n569_), .B1(new_n524_), .B2(new_n570_), .ZN(new_n1516_));
  OR2_X1    g1087(.A1(new_n1516_), .A2(KEYINPUT115), .ZN(new_n1517_));
  NAND2_X1  g1088(.A1(new_n1516_), .A2(KEYINPUT115), .ZN(new_n1518_));
  OAI211_X1 g1089(.A(new_n1517_), .B(new_n1518_), .C1(new_n537_), .C2(G273), .ZN(new_n1519_));
  NAND3_X1  g1090(.A1(new_n570_), .A2(G251), .A3(G411), .ZN(new_n1520_));
  NAND3_X1  g1091(.A1(G248), .A2(G273), .A3(G411), .ZN(new_n1521_));
  AND2_X1   g1092(.A1(new_n1521_), .A2(KEYINPUT116), .ZN(new_n1522_));
  NOR2_X1   g1093(.A1(new_n1521_), .A2(KEYINPUT116), .ZN(new_n1523_));
  OAI211_X1 g1094(.A(new_n1519_), .B(new_n1520_), .C1(new_n1522_), .C2(new_n1523_), .ZN(new_n1524_));
  NAND3_X1  g1095(.A1(G248), .A2(G281), .A3(G374), .ZN(new_n1525_));
  XNOR2_X1  g1096(.A(new_n1525_), .B(KEYINPUT117), .ZN(new_n1526_));
  NAND3_X1  g1097(.A1(new_n550_), .A2(G251), .A3(G374), .ZN(new_n1527_));
  AOI21_X1  g1098(.A(G374), .B1(new_n550_), .B2(G254), .ZN(new_n1528_));
  OAI21_X1  g1099(.A(new_n1528_), .B1(new_n524_), .B2(new_n550_), .ZN(new_n1529_));
  NAND3_X1  g1100(.A1(new_n1526_), .A2(new_n1527_), .A3(new_n1529_), .ZN(new_n1530_));
  XNOR2_X1  g1101(.A(new_n1524_), .B(new_n1530_), .ZN(new_n1531_));
  AOI21_X1  g1102(.A(G422), .B1(new_n611_), .B2(G254), .ZN(new_n1532_));
  OAI21_X1  g1103(.A(new_n1532_), .B1(new_n611_), .B2(new_n524_), .ZN(new_n1533_));
  OAI221_X1 g1104(.A(new_n1533_), .B1(new_n1359_), .B2(new_n615_), .C1(new_n544_), .C2(new_n614_), .ZN(new_n1534_));
  XOR2_X1   g1105(.A(new_n1531_), .B(new_n1534_), .Z(new_n1535_));
  AOI21_X1  g1106(.A(G4091), .B1(new_n1515_), .B2(new_n1535_), .ZN(new_n1536_));
  OAI21_X1  g1107(.A(new_n1536_), .B1(new_n1535_), .B2(new_n1515_), .ZN(new_n1537_));
  NOR2_X1   g1108(.A1(new_n1537_), .A2(G4092), .ZN(new_n1538_));
  XNOR2_X1  g1109(.A(new_n1538_), .B(KEYINPUT121), .ZN(new_n1539_));
  INV_X1    g1110(.A(new_n674_), .ZN(new_n1540_));
  INV_X1    g1111(.A(new_n821_), .ZN(new_n1541_));
  NAND4_X1  g1112(.A1(new_n973_), .A2(new_n969_), .A3(new_n972_), .A4(new_n1541_), .ZN(new_n1542_));
  AOI21_X1  g1113(.A(new_n683_), .B1(new_n985_), .B2(new_n665_), .ZN(new_n1543_));
  OAI21_X1  g1114(.A(new_n821_), .B1(new_n971_), .B2(new_n1543_), .ZN(new_n1544_));
  NAND2_X1  g1115(.A1(new_n1542_), .A2(new_n1544_), .ZN(new_n1545_));
  NAND2_X1  g1116(.A1(new_n1545_), .A2(KEYINPUT108), .ZN(new_n1546_));
  NAND2_X1  g1117(.A1(new_n954_), .A2(new_n953_), .ZN(new_n1547_));
  AND2_X1   g1118(.A1(new_n944_), .A2(new_n947_), .ZN(new_n1548_));
  NOR2_X1   g1119(.A1(new_n826_), .A2(new_n943_), .ZN(new_n1549_));
  NAND3_X1  g1120(.A1(new_n1547_), .A2(new_n1548_), .A3(new_n1549_), .ZN(new_n1550_));
  AND3_X1   g1121(.A1(new_n987_), .A2(new_n988_), .A3(new_n989_), .ZN(new_n1551_));
  NAND2_X1  g1122(.A1(new_n1550_), .A2(new_n1551_), .ZN(new_n1552_));
  INV_X1    g1123(.A(KEYINPUT108), .ZN(new_n1553_));
  NAND3_X1  g1124(.A1(new_n1542_), .A2(new_n1553_), .A3(new_n1544_), .ZN(new_n1554_));
  NAND4_X1  g1125(.A1(new_n1547_), .A2(new_n1548_), .A3(new_n1549_), .A4(new_n990_), .ZN(new_n1555_));
  AND4_X1   g1126(.A1(new_n1546_), .A2(new_n1552_), .A3(new_n1554_), .A4(new_n1555_), .ZN(new_n1556_));
  AOI22_X1  g1127(.A1(new_n1552_), .A2(new_n1555_), .B1(new_n1546_), .B2(new_n1554_), .ZN(new_n1557_));
  OAI21_X1  g1128(.A(new_n784_), .B1(new_n1556_), .B2(new_n1557_), .ZN(new_n1558_));
  AOI21_X1  g1129(.A(new_n990_), .B1(new_n955_), .B2(new_n1549_), .ZN(new_n1559_));
  INV_X1    g1130(.A(new_n1555_), .ZN(new_n1560_));
  INV_X1    g1131(.A(new_n1554_), .ZN(new_n1561_));
  AOI21_X1  g1132(.A(new_n1553_), .B1(new_n1542_), .B2(new_n1544_), .ZN(new_n1562_));
  OAI22_X1  g1133(.A1(new_n1559_), .A2(new_n1560_), .B1(new_n1561_), .B2(new_n1562_), .ZN(new_n1563_));
  NAND4_X1  g1134(.A1(new_n1552_), .A2(new_n1546_), .A3(new_n1554_), .A4(new_n1555_), .ZN(new_n1564_));
  NAND3_X1  g1135(.A1(new_n1563_), .A2(new_n785_), .A3(new_n1564_), .ZN(new_n1565_));
  NAND3_X1  g1136(.A1(new_n1558_), .A2(KEYINPUT109), .A3(new_n1565_), .ZN(new_n1566_));
  AOI21_X1  g1137(.A(new_n785_), .B1(new_n1563_), .B2(new_n1564_), .ZN(new_n1567_));
  INV_X1    g1138(.A(KEYINPUT109), .ZN(new_n1568_));
  NAND2_X1  g1139(.A1(new_n1567_), .A2(new_n1568_), .ZN(new_n1569_));
  AOI21_X1  g1140(.A(new_n1540_), .B1(new_n1566_), .B2(new_n1569_), .ZN(new_n1570_));
  AND3_X1   g1141(.A1(new_n1563_), .A2(new_n785_), .A3(new_n1564_), .ZN(new_n1571_));
  OAI21_X1  g1142(.A(new_n1540_), .B1(new_n1571_), .B2(new_n1567_), .ZN(new_n1572_));
  NAND2_X1  g1143(.A1(new_n1572_), .A2(KEYINPUT110), .ZN(new_n1573_));
  NOR2_X1   g1144(.A1(new_n1570_), .A2(new_n1573_), .ZN(new_n1574_));
  AOI211_X1 g1145(.A(KEYINPUT110), .B(new_n1540_), .C1(new_n1566_), .C2(new_n1569_), .ZN(new_n1575_));
  OAI21_X1  g1146(.A(new_n632_), .B1(new_n1574_), .B2(new_n1575_), .ZN(new_n1576_));
  NAND2_X1  g1147(.A1(new_n1566_), .A2(new_n1569_), .ZN(new_n1577_));
  INV_X1    g1148(.A(KEYINPUT110), .ZN(new_n1578_));
  NAND3_X1  g1149(.A1(new_n1577_), .A2(new_n1578_), .A3(new_n674_), .ZN(new_n1579_));
  OAI211_X1 g1150(.A(new_n1579_), .B(new_n783_), .C1(new_n1570_), .C2(new_n1573_), .ZN(new_n1580_));
  NAND2_X1  g1151(.A1(new_n1576_), .A2(new_n1580_), .ZN(new_n1581_));
  NAND2_X1  g1152(.A1(new_n1581_), .A2(new_n685_), .ZN(new_n1582_));
  AOI21_X1  g1153(.A(new_n674_), .B1(new_n1566_), .B2(new_n1569_), .ZN(new_n1583_));
  OAI21_X1  g1154(.A(new_n674_), .B1(new_n1571_), .B2(new_n1567_), .ZN(new_n1584_));
  NAND2_X1  g1155(.A1(new_n1584_), .A2(new_n783_), .ZN(new_n1585_));
  OAI21_X1  g1156(.A(new_n786_), .B1(new_n1583_), .B2(new_n1585_), .ZN(new_n1586_));
  OAI21_X1  g1157(.A(new_n1579_), .B1(new_n1570_), .B2(new_n1573_), .ZN(new_n1587_));
  AOI21_X1  g1158(.A(new_n1586_), .B1(new_n1587_), .B2(new_n632_), .ZN(new_n1588_));
  INV_X1    g1159(.A(new_n1588_), .ZN(new_n1589_));
  NAND3_X1  g1160(.A1(new_n1582_), .A2(new_n1589_), .A3(new_n828_), .ZN(new_n1590_));
  INV_X1    g1161(.A(G1497), .ZN(new_n1591_));
  AOI21_X1  g1162(.A(new_n684_), .B1(new_n1576_), .B2(new_n1580_), .ZN(new_n1592_));
  OAI21_X1  g1163(.A(new_n646_), .B1(new_n1592_), .B2(new_n1588_), .ZN(new_n1593_));
  NAND3_X1  g1164(.A1(new_n1590_), .A2(new_n1591_), .A3(new_n1593_), .ZN(new_n1594_));
  INV_X1    g1165(.A(new_n698_), .ZN(new_n1595_));
  OAI22_X1  g1166(.A1(new_n1043_), .A2(KEYINPUT99), .B1(new_n1595_), .B2(new_n693_), .ZN(new_n1596_));
  AOI21_X1  g1167(.A(new_n1596_), .B1(KEYINPUT99), .B2(new_n1043_), .ZN(new_n1597_));
  XNOR2_X1  g1168(.A(new_n1597_), .B(new_n1045_), .ZN(new_n1598_));
  XNOR2_X1  g1169(.A(new_n1598_), .B(new_n695_), .ZN(new_n1599_));
  OAI21_X1  g1170(.A(KEYINPUT100), .B1(new_n1598_), .B2(new_n1048_), .ZN(new_n1600_));
  XNOR2_X1  g1171(.A(new_n704_), .B(new_n700_), .ZN(new_n1601_));
  NAND2_X1  g1172(.A1(new_n1600_), .A2(new_n1601_), .ZN(new_n1602_));
  XNOR2_X1  g1173(.A(new_n1599_), .B(new_n1602_), .ZN(new_n1603_));
  OR3_X1    g1174(.A1(new_n1603_), .A2(KEYINPUT101), .A3(new_n711_), .ZN(new_n1604_));
  OAI21_X1  g1175(.A(KEYINPUT101), .B1(new_n1603_), .B2(new_n711_), .ZN(new_n1605_));
  OAI21_X1  g1176(.A(new_n834_), .B1(new_n688_), .B2(new_n1591_), .ZN(new_n1606_));
  INV_X1    g1177(.A(new_n1606_), .ZN(new_n1607_));
  AOI21_X1  g1178(.A(new_n1607_), .B1(new_n1603_), .B2(new_n711_), .ZN(new_n1608_));
  NAND3_X1  g1179(.A1(new_n1604_), .A2(new_n1605_), .A3(new_n1608_), .ZN(new_n1609_));
  NAND2_X1  g1180(.A1(new_n692_), .A2(new_n698_), .ZN(new_n1610_));
  NAND2_X1  g1181(.A1(new_n1610_), .A2(new_n813_), .ZN(new_n1611_));
  NAND2_X1  g1182(.A1(new_n1611_), .A2(KEYINPUT102), .ZN(new_n1612_));
  INV_X1    g1183(.A(KEYINPUT102), .ZN(new_n1613_));
  NAND3_X1  g1184(.A1(new_n1610_), .A2(new_n813_), .A3(new_n1613_), .ZN(new_n1614_));
  AND3_X1   g1185(.A1(new_n1612_), .A2(new_n816_), .A3(new_n1614_), .ZN(new_n1615_));
  AOI21_X1  g1186(.A(new_n816_), .B1(new_n1612_), .B2(new_n1614_), .ZN(new_n1616_));
  OAI21_X1  g1187(.A(new_n695_), .B1(new_n1615_), .B2(new_n1616_), .ZN(new_n1617_));
  NAND2_X1  g1188(.A1(new_n1612_), .A2(new_n1614_), .ZN(new_n1618_));
  INV_X1    g1189(.A(new_n816_), .ZN(new_n1619_));
  NAND2_X1  g1190(.A1(new_n1618_), .A2(new_n1619_), .ZN(new_n1620_));
  NAND3_X1  g1191(.A1(new_n1612_), .A2(new_n816_), .A3(new_n1614_), .ZN(new_n1621_));
  NAND3_X1  g1192(.A1(new_n1620_), .A2(new_n1048_), .A3(new_n1621_), .ZN(new_n1622_));
  NAND2_X1  g1193(.A1(new_n1617_), .A2(new_n1622_), .ZN(new_n1623_));
  AOI21_X1  g1194(.A(new_n701_), .B1(new_n1623_), .B2(KEYINPUT105), .ZN(new_n1624_));
  INV_X1    g1195(.A(KEYINPUT105), .ZN(new_n1625_));
  NAND3_X1  g1196(.A1(new_n1617_), .A2(new_n1622_), .A3(new_n1625_), .ZN(new_n1626_));
  AOI21_X1  g1197(.A(new_n811_), .B1(new_n1624_), .B2(new_n1626_), .ZN(new_n1627_));
  NAND3_X1  g1198(.A1(new_n1617_), .A2(new_n1622_), .A3(KEYINPUT103), .ZN(new_n1628_));
  INV_X1    g1199(.A(KEYINPUT103), .ZN(new_n1629_));
  OAI211_X1 g1200(.A(new_n1629_), .B(new_n695_), .C1(new_n1615_), .C2(new_n1616_), .ZN(new_n1630_));
  NAND2_X1  g1201(.A1(new_n1628_), .A2(new_n1630_), .ZN(new_n1631_));
  AOI21_X1  g1202(.A(KEYINPUT104), .B1(new_n1631_), .B2(new_n701_), .ZN(new_n1632_));
  INV_X1    g1203(.A(KEYINPUT104), .ZN(new_n1633_));
  AOI211_X1 g1204(.A(new_n1633_), .B(new_n700_), .C1(new_n1628_), .C2(new_n1630_), .ZN(new_n1634_));
  OAI21_X1  g1205(.A(new_n1627_), .B1(new_n1632_), .B2(new_n1634_), .ZN(new_n1635_));
  INV_X1    g1206(.A(KEYINPUT106), .ZN(new_n1636_));
  NAND2_X1  g1207(.A1(new_n1635_), .A2(new_n1636_), .ZN(new_n1637_));
  OAI211_X1 g1208(.A(new_n1627_), .B(KEYINPUT106), .C1(new_n1632_), .C2(new_n1634_), .ZN(new_n1638_));
  OAI22_X1  g1209(.A1(new_n1632_), .A2(new_n1634_), .B1(new_n701_), .B2(new_n1631_), .ZN(new_n1639_));
  AOI22_X1  g1210(.A1(new_n1637_), .A2(new_n1638_), .B1(new_n811_), .B2(new_n1639_), .ZN(new_n1640_));
  OAI21_X1  g1211(.A(new_n1607_), .B1(new_n1640_), .B2(new_n711_), .ZN(new_n1641_));
  NAND2_X1  g1212(.A1(new_n1637_), .A2(new_n1638_), .ZN(new_n1642_));
  NAND2_X1  g1213(.A1(new_n1639_), .A2(new_n811_), .ZN(new_n1643_));
  AND3_X1   g1214(.A1(new_n1642_), .A2(new_n711_), .A3(new_n1643_), .ZN(new_n1644_));
  OAI21_X1  g1215(.A(new_n1609_), .B1(new_n1641_), .B2(new_n1644_), .ZN(new_n1645_));
  NAND2_X1  g1216(.A1(new_n787_), .A2(new_n663_), .ZN(new_n1646_));
  NAND2_X1  g1217(.A1(new_n1646_), .A2(new_n972_), .ZN(new_n1647_));
  NAND2_X1  g1218(.A1(new_n971_), .A2(new_n663_), .ZN(new_n1648_));
  INV_X1    g1219(.A(new_n675_), .ZN(new_n1649_));
  OAI211_X1 g1220(.A(new_n1647_), .B(new_n1648_), .C1(new_n1649_), .C2(new_n990_), .ZN(new_n1650_));
  INV_X1    g1221(.A(new_n1648_), .ZN(new_n1651_));
  AOI21_X1  g1222(.A(new_n971_), .B1(new_n787_), .B2(new_n663_), .ZN(new_n1652_));
  OAI211_X1 g1223(.A(new_n675_), .B(new_n1551_), .C1(new_n1651_), .C2(new_n1652_), .ZN(new_n1653_));
  INV_X1    g1224(.A(KEYINPUT107), .ZN(new_n1654_));
  NAND3_X1  g1225(.A1(new_n1650_), .A2(new_n1653_), .A3(new_n1654_), .ZN(new_n1655_));
  INV_X1    g1226(.A(new_n789_), .ZN(new_n1656_));
  NOR2_X1   g1227(.A1(new_n1550_), .A2(new_n1656_), .ZN(new_n1657_));
  NAND2_X1  g1228(.A1(new_n1551_), .A2(new_n675_), .ZN(new_n1658_));
  NAND4_X1  g1229(.A1(new_n1658_), .A2(KEYINPUT107), .A3(new_n1647_), .A4(new_n1648_), .ZN(new_n1659_));
  NAND3_X1  g1230(.A1(new_n1655_), .A2(new_n1657_), .A3(new_n1659_), .ZN(new_n1660_));
  NAND3_X1  g1231(.A1(new_n955_), .A2(new_n789_), .A3(new_n1549_), .ZN(new_n1661_));
  NAND3_X1  g1232(.A1(new_n1661_), .A2(new_n1650_), .A3(new_n1653_), .ZN(new_n1662_));
  NAND2_X1  g1233(.A1(new_n1660_), .A2(new_n1662_), .ZN(new_n1663_));
  NAND2_X1  g1234(.A1(new_n1663_), .A2(new_n784_), .ZN(new_n1664_));
  NAND3_X1  g1235(.A1(new_n1660_), .A2(new_n785_), .A3(new_n1662_), .ZN(new_n1665_));
  AOI21_X1  g1236(.A(new_n674_), .B1(new_n1664_), .B2(new_n1665_), .ZN(new_n1666_));
  NAND3_X1  g1237(.A1(new_n1655_), .A2(new_n1661_), .A3(new_n1659_), .ZN(new_n1667_));
  NAND4_X1  g1238(.A1(new_n1650_), .A2(new_n1653_), .A3(new_n955_), .A4(new_n1549_), .ZN(new_n1668_));
  NAND3_X1  g1239(.A1(new_n1667_), .A2(new_n784_), .A3(new_n1668_), .ZN(new_n1669_));
  AND3_X1   g1240(.A1(new_n1665_), .A2(new_n1669_), .A3(new_n674_), .ZN(new_n1670_));
  NOR3_X1   g1241(.A1(new_n1666_), .A2(new_n1670_), .A3(new_n783_), .ZN(new_n1671_));
  INV_X1    g1242(.A(new_n1665_), .ZN(new_n1672_));
  AOI21_X1  g1243(.A(new_n785_), .B1(new_n1660_), .B2(new_n1662_), .ZN(new_n1673_));
  OAI21_X1  g1244(.A(new_n1540_), .B1(new_n1672_), .B2(new_n1673_), .ZN(new_n1674_));
  NAND3_X1  g1245(.A1(new_n1665_), .A2(new_n1669_), .A3(new_n674_), .ZN(new_n1675_));
  AOI21_X1  g1246(.A(new_n632_), .B1(new_n1674_), .B2(new_n1675_), .ZN(new_n1676_));
  OAI21_X1  g1247(.A(new_n685_), .B1(new_n1671_), .B2(new_n1676_), .ZN(new_n1677_));
  NAND3_X1  g1248(.A1(new_n1674_), .A2(new_n632_), .A3(new_n1675_), .ZN(new_n1678_));
  OAI21_X1  g1249(.A(new_n674_), .B1(new_n1672_), .B2(new_n1673_), .ZN(new_n1679_));
  NAND3_X1  g1250(.A1(new_n1665_), .A2(new_n1669_), .A3(new_n1540_), .ZN(new_n1680_));
  NAND3_X1  g1251(.A1(new_n1679_), .A2(new_n783_), .A3(new_n1680_), .ZN(new_n1681_));
  NAND3_X1  g1252(.A1(new_n1678_), .A2(new_n1681_), .A3(new_n786_), .ZN(new_n1682_));
  NAND3_X1  g1253(.A1(new_n1677_), .A2(new_n1682_), .A3(new_n828_), .ZN(new_n1683_));
  NAND2_X1  g1254(.A1(new_n1683_), .A2(KEYINPUT112), .ZN(new_n1684_));
  INV_X1    g1255(.A(KEYINPUT112), .ZN(new_n1685_));
  NAND4_X1  g1256(.A1(new_n1677_), .A2(new_n1682_), .A3(new_n1685_), .A4(new_n828_), .ZN(new_n1686_));
  NAND2_X1  g1257(.A1(new_n1677_), .A2(new_n1682_), .ZN(new_n1687_));
  NAND2_X1  g1258(.A1(new_n1687_), .A2(new_n646_), .ZN(new_n1688_));
  NAND3_X1  g1259(.A1(new_n1684_), .A2(new_n1686_), .A3(new_n1688_), .ZN(new_n1689_));
  AOI21_X1  g1260(.A(new_n1645_), .B1(new_n1689_), .B2(G1497), .ZN(new_n1690_));
  NAND2_X1  g1261(.A1(new_n1594_), .A2(new_n1690_), .ZN(new_n1691_));
  INV_X1    g1262(.A(KEYINPUT113), .ZN(new_n1692_));
  NAND2_X1  g1263(.A1(new_n1691_), .A2(new_n1692_), .ZN(new_n1693_));
  NAND3_X1  g1264(.A1(new_n1594_), .A2(new_n1690_), .A3(KEYINPUT113), .ZN(new_n1694_));
  NAND2_X1  g1265(.A1(new_n1693_), .A2(new_n1694_), .ZN(new_n1695_));
  INV_X1    g1266(.A(new_n1645_), .ZN(new_n1696_));
  NAND2_X1  g1267(.A1(new_n1590_), .A2(KEYINPUT111), .ZN(new_n1697_));
  INV_X1    g1268(.A(KEYINPUT111), .ZN(new_n1698_));
  NAND4_X1  g1269(.A1(new_n1582_), .A2(new_n1589_), .A3(new_n1698_), .A4(new_n828_), .ZN(new_n1699_));
  NAND4_X1  g1270(.A1(new_n1697_), .A2(new_n1591_), .A3(new_n1699_), .A4(new_n1593_), .ZN(new_n1700_));
  INV_X1    g1271(.A(new_n1683_), .ZN(new_n1701_));
  NAND2_X1  g1272(.A1(new_n1678_), .A2(new_n1681_), .ZN(new_n1702_));
  NAND2_X1  g1273(.A1(new_n1702_), .A2(new_n950_), .ZN(new_n1703_));
  OAI21_X1  g1274(.A(new_n783_), .B1(new_n1666_), .B2(new_n1670_), .ZN(new_n1704_));
  NAND3_X1  g1275(.A1(new_n1704_), .A2(new_n1678_), .A3(new_n684_), .ZN(new_n1705_));
  AOI21_X1  g1276(.A(new_n647_), .B1(new_n1703_), .B2(new_n1705_), .ZN(new_n1706_));
  OAI21_X1  g1277(.A(G1497), .B1(new_n1701_), .B2(new_n1706_), .ZN(new_n1707_));
  AOI21_X1  g1278(.A(new_n1696_), .B1(new_n1700_), .B2(new_n1707_), .ZN(new_n1708_));
  OAI21_X1  g1279(.A(G4091), .B1(new_n1695_), .B2(new_n1708_), .ZN(new_n1709_));
  OAI211_X1 g1280(.A(new_n1483_), .B(new_n1539_), .C1(new_n1709_), .C2(G4092), .ZN(G882));
  OAI21_X1  g1281(.A(G4087), .B1(G14), .B2(G4088), .ZN(new_n1711_));
  INV_X1    g1282(.A(G64), .ZN(new_n1712_));
  AOI21_X1  g1283(.A(new_n1711_), .B1(new_n1712_), .B2(G4088), .ZN(new_n1713_));
  AOI21_X1  g1284(.A(G4092), .B1(new_n1371_), .B2(new_n861_), .ZN(new_n1714_));
  INV_X1    g1285(.A(new_n1714_), .ZN(new_n1715_));
  AOI21_X1  g1286(.A(new_n1715_), .B1(new_n1480_), .B2(G4091), .ZN(new_n1716_));
  NAND2_X1  g1287(.A1(G94), .A2(G4092), .ZN(new_n1717_));
  XOR2_X1   g1288(.A(new_n1717_), .B(KEYINPUT123), .Z(new_n1718_));
  INV_X1    g1289(.A(new_n1718_), .ZN(new_n1719_));
  OAI211_X1 g1290(.A(KEYINPUT124), .B(new_n1106_), .C1(new_n1716_), .C2(new_n1719_), .ZN(new_n1720_));
  INV_X1    g1291(.A(KEYINPUT124), .ZN(new_n1721_));
  AOI21_X1  g1292(.A(new_n1471_), .B1(new_n1460_), .B2(new_n736_), .ZN(new_n1722_));
  AOI21_X1  g1293(.A(new_n1477_), .B1(new_n1466_), .B2(new_n1722_), .ZN(new_n1723_));
  NAND2_X1  g1294(.A1(new_n1461_), .A2(new_n1462_), .ZN(new_n1724_));
  OAI21_X1  g1295(.A(new_n1417_), .B1(new_n1723_), .B2(new_n1724_), .ZN(new_n1725_));
  NAND2_X1  g1296(.A1(new_n1725_), .A2(new_n1398_), .ZN(new_n1726_));
  NAND3_X1  g1297(.A1(new_n1478_), .A2(new_n1417_), .A3(new_n1475_), .ZN(new_n1727_));
  NAND3_X1  g1298(.A1(new_n1726_), .A2(G4091), .A3(new_n1727_), .ZN(new_n1728_));
  AOI21_X1  g1299(.A(new_n1719_), .B1(new_n1728_), .B2(new_n1714_), .ZN(new_n1729_));
  OAI21_X1  g1300(.A(new_n1721_), .B1(new_n1729_), .B2(new_n1107_), .ZN(new_n1730_));
  AOI21_X1  g1301(.A(new_n1713_), .B1(new_n1720_), .B2(new_n1730_), .ZN(new_n1731_));
  NAND2_X1  g1302(.A1(G97), .A2(G4092), .ZN(new_n1732_));
  INV_X1    g1303(.A(new_n1732_), .ZN(new_n1733_));
  NAND2_X1  g1304(.A1(new_n1537_), .A2(new_n854_), .ZN(new_n1734_));
  INV_X1    g1305(.A(new_n1734_), .ZN(new_n1735_));
  AOI21_X1  g1306(.A(new_n1733_), .B1(new_n1709_), .B2(new_n1735_), .ZN(new_n1736_));
  INV_X1    g1307(.A(KEYINPUT122), .ZN(new_n1737_));
  NOR3_X1   g1308(.A1(new_n1736_), .A2(new_n1737_), .A3(new_n904_), .ZN(new_n1738_));
  AND3_X1   g1309(.A1(new_n1594_), .A2(new_n1690_), .A3(KEYINPUT113), .ZN(new_n1739_));
  AOI21_X1  g1310(.A(KEYINPUT113), .B1(new_n1594_), .B2(new_n1690_), .ZN(new_n1740_));
  NOR2_X1   g1311(.A1(new_n1739_), .A2(new_n1740_), .ZN(new_n1741_));
  NOR3_X1   g1312(.A1(new_n1592_), .A2(new_n646_), .A3(new_n1588_), .ZN(new_n1742_));
  OAI211_X1 g1313(.A(new_n1591_), .B(new_n1593_), .C1(new_n1742_), .C2(new_n1698_), .ZN(new_n1743_));
  INV_X1    g1314(.A(new_n1699_), .ZN(new_n1744_));
  OAI21_X1  g1315(.A(new_n1707_), .B1(new_n1743_), .B2(new_n1744_), .ZN(new_n1745_));
  NAND2_X1  g1316(.A1(new_n1745_), .A2(new_n1645_), .ZN(new_n1746_));
  AOI21_X1  g1317(.A(new_n861_), .B1(new_n1741_), .B2(new_n1746_), .ZN(new_n1747_));
  OAI21_X1  g1318(.A(new_n1732_), .B1(new_n1747_), .B2(new_n1734_), .ZN(new_n1748_));
  AOI21_X1  g1319(.A(KEYINPUT122), .B1(new_n1748_), .B2(new_n903_), .ZN(new_n1749_));
  OAI21_X1  g1320(.A(new_n1731_), .B1(new_n1738_), .B2(new_n1749_), .ZN(G767));
  NAND2_X1  g1321(.A1(new_n1712_), .A2(G4089), .ZN(new_n1751_));
  OAI211_X1 g1322(.A(new_n1751_), .B(G4090), .C1(G14), .C2(G4089), .ZN(new_n1752_));
  NAND2_X1  g1323(.A1(new_n1728_), .A2(new_n1714_), .ZN(new_n1753_));
  NAND2_X1  g1324(.A1(new_n1753_), .A2(new_n1718_), .ZN(new_n1754_));
  AOI21_X1  g1325(.A(KEYINPUT125), .B1(new_n1754_), .B2(new_n1122_), .ZN(new_n1755_));
  INV_X1    g1326(.A(KEYINPUT125), .ZN(new_n1756_));
  NOR3_X1   g1327(.A1(new_n1729_), .A2(new_n1756_), .A3(new_n1134_), .ZN(new_n1757_));
  OAI221_X1 g1328(.A(new_n1752_), .B1(new_n1736_), .B2(new_n941_), .C1(new_n1755_), .C2(new_n1757_), .ZN(G807));
  NAND3_X1  g1329(.A1(new_n1081_), .A2(G176), .A3(G1690), .ZN(new_n1759_));
  OR2_X1    g1330(.A1(new_n1759_), .A2(KEYINPUT126), .ZN(new_n1760_));
  NAND3_X1  g1331(.A1(G179), .A2(G1689), .A3(G1690), .ZN(new_n1761_));
  NAND2_X1  g1332(.A1(new_n1759_), .A2(KEYINPUT126), .ZN(new_n1762_));
  NAND3_X1  g1333(.A1(new_n1760_), .A2(new_n1761_), .A3(new_n1762_), .ZN(new_n1763_));
  AOI21_X1  g1334(.A(new_n1763_), .B1(new_n1754_), .B2(new_n1089_), .ZN(new_n1764_));
  OAI21_X1  g1335(.A(new_n1764_), .B1(new_n1083_), .B2(new_n1736_), .ZN(new_n1765_));
  NAND2_X1  g1336(.A1(new_n1765_), .A2(G137), .ZN(G658));
  NAND3_X1  g1337(.A1(new_n1096_), .A2(G176), .A3(G1694), .ZN(new_n1767_));
  INV_X1    g1338(.A(KEYINPUT127), .ZN(new_n1768_));
  OR2_X1    g1339(.A1(new_n1767_), .A2(new_n1768_), .ZN(new_n1769_));
  NAND3_X1  g1340(.A1(G179), .A2(G1691), .A3(G1694), .ZN(new_n1770_));
  NAND2_X1  g1341(.A1(new_n1767_), .A2(new_n1768_), .ZN(new_n1771_));
  NAND3_X1  g1342(.A1(new_n1769_), .A2(new_n1770_), .A3(new_n1771_), .ZN(new_n1772_));
  AOI21_X1  g1343(.A(new_n1772_), .B1(new_n1754_), .B2(new_n1176_), .ZN(new_n1773_));
  OAI21_X1  g1344(.A(new_n1773_), .B1(new_n1179_), .B2(new_n1736_), .ZN(new_n1774_));
  NAND2_X1  g1345(.A1(new_n1774_), .A2(G137), .ZN(G690));
endmodule


