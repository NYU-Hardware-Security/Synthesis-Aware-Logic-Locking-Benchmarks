//Secret key is'1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_c1908" written by ABC on Sun Nov 20 19:50:24 2022

module locked_c1908 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64, KEYINPUT65,
    KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70, KEYINPUT71,
    KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76, KEYINPUT77,
    KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82, KEYINPUT83,
    KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88, KEYINPUT89,
    KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94, KEYINPUT95,
    KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99, KEYINPUT100,
    KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104, KEYINPUT105,
    KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109, KEYINPUT110,
    KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114, KEYINPUT115,
    KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119, KEYINPUT120,
    KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124, KEYINPUT125,
    KEYINPUT126, KEYINPUT127, G101, G104, G107, G110, G113, G116, G119,
    G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217,
    G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902,
    G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, KEYINPUT64,
    KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69, KEYINPUT70,
    KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75, KEYINPUT76,
    KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81, KEYINPUT82,
    KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87, KEYINPUT88,
    KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93, KEYINPUT94,
    KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, G101, G104, G107, G110, G113,
    G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210,
    G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898,
    G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_;
  INV_X1    g000(.A(G469), .ZN(new_n187_));
  XNOR2_X1  g001(.A(KEYINPUT0), .B(G902), .ZN(new_n188_));
  INV_X1    g002(.A(G131), .ZN(new_n189_));
  INV_X1    g003(.A(G134), .ZN(new_n190_));
  NAND2_X1  g004(.A1(new_n190_), .A2(G137), .ZN(new_n191_));
  INV_X1    g005(.A(G137), .ZN(new_n192_));
  AND3_X1   g006(.A1(new_n192_), .A2(KEYINPUT27), .A3(G134), .ZN(new_n193_));
  AOI21_X1  g007(.A(KEYINPUT27), .B1(new_n192_), .B2(G134), .ZN(new_n194_));
  OAI211_X1 g008(.A(new_n189_), .B(new_n191_), .C1(new_n193_), .C2(new_n194_), .ZN(new_n195_));
  NAND2_X1  g009(.A1(new_n195_), .A2(KEYINPUT28), .ZN(new_n196_));
  NAND2_X1  g010(.A1(new_n192_), .A2(G134), .ZN(new_n197_));
  INV_X1    g011(.A(KEYINPUT27), .ZN(new_n198_));
  NAND2_X1  g012(.A1(new_n197_), .A2(new_n198_), .ZN(new_n199_));
  NAND3_X1  g013(.A1(new_n192_), .A2(KEYINPUT27), .A3(G134), .ZN(new_n200_));
  NAND2_X1  g014(.A1(new_n199_), .A2(new_n200_), .ZN(new_n201_));
  INV_X1    g015(.A(KEYINPUT28), .ZN(new_n202_));
  NAND4_X1  g016(.A1(new_n201_), .A2(new_n202_), .A3(new_n189_), .A4(new_n191_), .ZN(new_n203_));
  OAI21_X1  g017(.A(new_n191_), .B1(new_n193_), .B2(new_n194_), .ZN(new_n204_));
  NAND2_X1  g018(.A1(new_n204_), .A2(G131), .ZN(new_n205_));
  NAND3_X1  g019(.A1(new_n196_), .A2(new_n203_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g020(.A(G104), .ZN(new_n207_));
  NAND2_X1  g021(.A1(new_n207_), .A2(KEYINPUT7), .ZN(new_n208_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n209_));
  NAND2_X1  g023(.A1(new_n209_), .A2(G104), .ZN(new_n210_));
  INV_X1    g024(.A(G107), .ZN(new_n211_));
  NAND3_X1  g025(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g026(.A(KEYINPUT10), .ZN(new_n213_));
  NAND2_X1  g027(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g028(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT10), .A4(new_n211_), .ZN(new_n215_));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216_));
  AOI21_X1  g030(.A(new_n216_), .B1(new_n207_), .B2(G107), .ZN(new_n217_));
  NOR3_X1   g031(.A1(new_n211_), .A2(KEYINPUT11), .A3(G104), .ZN(new_n218_));
  NOR2_X1   g032(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g033(.A1(new_n214_), .A2(new_n215_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g034(.A1(new_n220_), .A2(G101), .ZN(new_n221_));
  NAND2_X1  g035(.A1(new_n221_), .A2(KEYINPUT12), .ZN(new_n222_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n223_));
  NAND3_X1  g037(.A1(new_n220_), .A2(new_n223_), .A3(G101), .ZN(new_n224_));
  NAND3_X1  g038(.A1(new_n211_), .A2(KEYINPUT6), .A3(G104), .ZN(new_n225_));
  INV_X1    g039(.A(KEYINPUT6), .ZN(new_n226_));
  OAI21_X1  g040(.A(new_n226_), .B1(new_n207_), .B2(G107), .ZN(new_n227_));
  XNOR2_X1  g041(.A(KEYINPUT7), .B(G104), .ZN(new_n228_));
  OAI211_X1 g042(.A(new_n225_), .B(new_n227_), .C1(new_n228_), .C2(new_n211_), .ZN(new_n229_));
  OAI21_X1  g043(.A(KEYINPUT9), .B1(new_n229_), .B2(G101), .ZN(new_n230_));
  NAND2_X1  g044(.A1(new_n208_), .A2(new_n210_), .ZN(new_n231_));
  NAND2_X1  g045(.A1(new_n231_), .A2(G107), .ZN(new_n232_));
  AND2_X1   g046(.A1(new_n227_), .A2(new_n225_), .ZN(new_n233_));
  INV_X1    g047(.A(KEYINPUT9), .ZN(new_n234_));
  INV_X1    g048(.A(G101), .ZN(new_n235_));
  NAND4_X1  g049(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  AOI22_X1  g050(.A1(new_n222_), .A2(new_n224_), .B1(new_n230_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g051(.A(G128), .ZN(new_n238_));
  INV_X1    g052(.A(G146), .ZN(new_n239_));
  NAND2_X1  g053(.A1(new_n239_), .A2(G143), .ZN(new_n240_));
  INV_X1    g054(.A(G143), .ZN(new_n241_));
  NAND2_X1  g055(.A1(new_n241_), .A2(G146), .ZN(new_n242_));
  AOI21_X1  g056(.A(new_n238_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244_));
  NAND3_X1  g058(.A1(new_n244_), .A2(new_n239_), .A3(G143), .ZN(new_n245_));
  AOI21_X1  g059(.A(KEYINPUT1), .B1(new_n241_), .B2(G146), .ZN(new_n246_));
  NOR2_X1   g060(.A1(new_n241_), .A2(G146), .ZN(new_n247_));
  OAI211_X1 g061(.A(new_n238_), .B(new_n245_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n249_));
  NAND2_X1  g063(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g064(.A(new_n244_), .B1(new_n239_), .B2(G143), .ZN(new_n251_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n240_), .ZN(new_n252_));
  NAND4_X1  g066(.A1(new_n252_), .A2(KEYINPUT2), .A3(new_n238_), .A4(new_n245_), .ZN(new_n253_));
  AOI21_X1  g067(.A(new_n243_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g068(.A1(new_n237_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g069(.A1(new_n230_), .A2(new_n236_), .ZN(new_n256_));
  AND3_X1   g070(.A1(new_n220_), .A2(new_n223_), .A3(G101), .ZN(new_n257_));
  AOI21_X1  g071(.A(new_n223_), .B1(new_n220_), .B2(G101), .ZN(new_n258_));
  OAI211_X1 g072(.A(new_n254_), .B(new_n256_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  INV_X1    g073(.A(new_n259_), .ZN(new_n260_));
  OAI21_X1  g074(.A(new_n206_), .B1(new_n255_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g075(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g076(.A(KEYINPUT26), .ZN(new_n263_));
  NAND2_X1  g077(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g078(.A1(new_n222_), .A2(new_n224_), .ZN(new_n265_));
  NAND4_X1  g079(.A1(new_n265_), .A2(KEYINPUT26), .A3(new_n254_), .A4(new_n256_), .ZN(new_n266_));
  INV_X1    g080(.A(new_n206_), .ZN(new_n267_));
  XNOR2_X1  g081(.A(new_n229_), .B(G101), .ZN(new_n268_));
  NAND2_X1  g082(.A1(new_n252_), .A2(new_n245_), .ZN(new_n269_));
  NAND2_X1  g083(.A1(new_n269_), .A2(G128), .ZN(new_n270_));
  NAND2_X1  g084(.A1(new_n270_), .A2(new_n248_), .ZN(new_n271_));
  NAND2_X1  g085(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g086(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .A4(new_n272_), .ZN(new_n273_));
  OR2_X1    g087(.A1(new_n273_), .A2(KEYINPUT30), .ZN(new_n274_));
  NAND2_X1  g088(.A1(new_n273_), .A2(KEYINPUT30), .ZN(new_n275_));
  AOI21_X1  g089(.A(new_n262_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g090(.A(G953), .ZN(new_n277_));
  NAND2_X1  g091(.A1(new_n277_), .A2(KEYINPUT25), .ZN(new_n278_));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n279_));
  NAND2_X1  g093(.A1(new_n279_), .A2(G953), .ZN(new_n280_));
  NAND2_X1  g094(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g095(.A1(new_n281_), .A2(G227), .ZN(new_n282_));
  XOR2_X1   g096(.A(G110), .B(G140), .Z(new_n283_));
  XOR2_X1   g097(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  INV_X1    g098(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g099(.A(new_n188_), .B1(new_n276_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g100(.A(new_n272_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n287_));
  INV_X1    g101(.A(new_n287_), .ZN(new_n288_));
  NAND4_X1  g102(.A1(new_n288_), .A2(KEYINPUT29), .A3(new_n267_), .A4(new_n264_), .ZN(new_n289_));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290_));
  NAND2_X1  g104(.A1(new_n273_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g105(.A(new_n264_), .ZN(new_n292_));
  OAI21_X1  g106(.A(new_n206_), .B1(new_n292_), .B2(new_n287_), .ZN(new_n293_));
  NAND3_X1  g107(.A1(new_n289_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g108(.A1(new_n294_), .A2(new_n284_), .ZN(new_n295_));
  AOI21_X1  g109(.A(new_n187_), .B1(new_n286_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g110(.A1(new_n294_), .A2(new_n285_), .ZN(new_n297_));
  AND2_X1   g111(.A1(new_n273_), .A2(KEYINPUT30), .ZN(new_n298_));
  NOR2_X1   g112(.A1(new_n273_), .A2(KEYINPUT30), .ZN(new_n299_));
  OAI211_X1 g113(.A(new_n284_), .B(new_n261_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  AND3_X1   g114(.A1(new_n297_), .A2(new_n300_), .A3(KEYINPUT31), .ZN(new_n301_));
  AOI21_X1  g115(.A(KEYINPUT31), .B1(new_n297_), .B2(new_n300_), .ZN(new_n302_));
  NOR2_X1   g116(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g117(.A1(new_n188_), .A2(G469), .ZN(new_n304_));
  AOI21_X1  g118(.A(new_n296_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g119(.A(G234), .ZN(new_n306_));
  OAI21_X1  g120(.A(G221), .B1(new_n306_), .B2(G902), .ZN(new_n307_));
  INV_X1    g121(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g122(.A(KEYINPUT32), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g123(.A1(new_n286_), .A2(new_n295_), .ZN(new_n310_));
  NAND2_X1  g124(.A1(new_n310_), .A2(G469), .ZN(new_n311_));
  NAND2_X1  g125(.A1(new_n297_), .A2(new_n300_), .ZN(new_n312_));
  INV_X1    g126(.A(KEYINPUT31), .ZN(new_n313_));
  NAND2_X1  g127(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g128(.A1(new_n297_), .A2(new_n300_), .A3(KEYINPUT31), .ZN(new_n315_));
  NAND3_X1  g129(.A1(new_n314_), .A2(new_n315_), .A3(new_n304_), .ZN(new_n316_));
  NAND2_X1  g130(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g131(.A(KEYINPUT32), .ZN(new_n318_));
  NAND3_X1  g132(.A1(new_n317_), .A2(new_n318_), .A3(new_n307_), .ZN(new_n319_));
  NAND2_X1  g133(.A1(new_n309_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g134(.A(G475), .ZN(new_n321_));
  OR2_X1    g135(.A1(KEYINPUT40), .A2(G237), .ZN(new_n322_));
  NAND2_X1  g136(.A1(KEYINPUT40), .A2(G237), .ZN(new_n323_));
  AOI22_X1  g137(.A1(new_n278_), .A2(new_n280_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g138(.A(G143), .B1(new_n324_), .B2(G214), .ZN(new_n325_));
  NAND2_X1  g139(.A1(new_n322_), .A2(new_n323_), .ZN(new_n326_));
  NAND4_X1  g140(.A1(new_n326_), .A2(new_n281_), .A3(G143), .A4(G214), .ZN(new_n327_));
  NAND2_X1  g141(.A1(new_n327_), .A2(KEYINPUT41), .ZN(new_n328_));
  INV_X1    g142(.A(KEYINPUT41), .ZN(new_n329_));
  NAND4_X1  g143(.A1(new_n324_), .A2(new_n329_), .A3(G143), .A4(G214), .ZN(new_n330_));
  AOI21_X1  g144(.A(new_n325_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g145(.A1(new_n331_), .A2(new_n189_), .ZN(new_n332_));
  NAND2_X1  g146(.A1(new_n328_), .A2(new_n330_), .ZN(new_n333_));
  INV_X1    g147(.A(G237), .ZN(new_n334_));
  NAND3_X1  g148(.A1(new_n334_), .A2(new_n277_), .A3(G214), .ZN(new_n335_));
  AOI21_X1  g149(.A(G131), .B1(new_n335_), .B2(new_n241_), .ZN(new_n336_));
  NAND2_X1  g150(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g151(.A(KEYINPUT42), .ZN(new_n338_));
  NAND2_X1  g152(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g153(.A1(new_n333_), .A2(KEYINPUT42), .A3(new_n336_), .ZN(new_n340_));
  AOI21_X1  g154(.A(new_n332_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g155(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343_));
  OR2_X1    g157(.A1(new_n343_), .A2(new_n239_), .ZN(new_n344_));
  NAND2_X1  g158(.A1(new_n343_), .A2(new_n239_), .ZN(new_n345_));
  NAND2_X1  g159(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g160(.A(new_n346_), .B(KEYINPUT39), .ZN(new_n347_));
  NAND2_X1  g161(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g162(.A(new_n346_), .ZN(new_n349_));
  AOI21_X1  g163(.A(new_n349_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n350_));
  OR2_X1    g164(.A1(new_n335_), .A2(KEYINPUT43), .ZN(new_n351_));
  AOI21_X1  g165(.A(G143), .B1(new_n335_), .B2(KEYINPUT43), .ZN(new_n352_));
  AOI22_X1  g166(.A1(new_n328_), .A2(new_n330_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g167(.A(new_n189_), .B1(new_n353_), .B2(KEYINPUT44), .ZN(new_n354_));
  NAND2_X1  g168(.A1(new_n351_), .A2(new_n352_), .ZN(new_n355_));
  NAND2_X1  g169(.A1(new_n333_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g170(.A(KEYINPUT44), .ZN(new_n357_));
  NAND2_X1  g171(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g172(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  AND3_X1   g173(.A1(new_n350_), .A2(KEYINPUT45), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g174(.A(KEYINPUT45), .B1(new_n350_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g175(.A(new_n348_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g176(.A(G113), .B(G122), .ZN(new_n363_));
  XNOR2_X1  g177(.A(new_n231_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g178(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g179(.A1(new_n362_), .A2(KEYINPUT47), .A3(new_n365_), .ZN(new_n366_));
  OAI211_X1 g180(.A(new_n348_), .B(new_n364_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n367_));
  NAND2_X1  g181(.A1(new_n367_), .A2(KEYINPUT46), .ZN(new_n368_));
  AOI21_X1  g182(.A(KEYINPUT46), .B1(new_n365_), .B2(KEYINPUT47), .ZN(new_n369_));
  OAI211_X1 g183(.A(new_n348_), .B(new_n369_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n370_));
  NAND3_X1  g184(.A1(new_n366_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g185(.A(G902), .ZN(new_n372_));
  NAND2_X1  g186(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g187(.A(new_n321_), .B1(new_n373_), .B2(KEYINPUT48), .ZN(new_n374_));
  INV_X1    g188(.A(KEYINPUT48), .ZN(new_n375_));
  NAND3_X1  g189(.A1(new_n371_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n376_));
  NAND3_X1  g190(.A1(new_n342_), .A2(KEYINPUT49), .A3(new_n349_), .ZN(new_n377_));
  INV_X1    g191(.A(KEYINPUT49), .ZN(new_n378_));
  OAI21_X1  g192(.A(new_n378_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n379_));
  NAND2_X1  g193(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g194(.A1(new_n360_), .A2(new_n361_), .ZN(new_n381_));
  OAI21_X1  g195(.A(new_n365_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g196(.A1(new_n382_), .A2(new_n367_), .ZN(new_n383_));
  NOR2_X1   g197(.A1(new_n188_), .A2(G475), .ZN(new_n384_));
  AOI22_X1  g198(.A1(new_n374_), .A2(new_n376_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g199(.A(new_n385_), .ZN(new_n386_));
  OAI211_X1 g200(.A(new_n281_), .B(G952), .C1(new_n306_), .C2(new_n334_), .ZN(new_n387_));
  XNOR2_X1  g201(.A(new_n387_), .B(KEYINPUT50), .ZN(new_n388_));
  AOI21_X1  g202(.A(new_n372_), .B1(G234), .B2(G237), .ZN(new_n389_));
  INV_X1    g203(.A(G898), .ZN(new_n390_));
  AND3_X1   g204(.A1(new_n389_), .A2(new_n390_), .A3(G953), .ZN(new_n391_));
  OR2_X1    g205(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g206(.A(new_n392_), .B(KEYINPUT51), .Z(new_n393_));
  INV_X1    g207(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g208(.A(G478), .ZN(new_n395_));
  INV_X1    g209(.A(new_n188_), .ZN(new_n396_));
  INV_X1    g210(.A(G116), .ZN(new_n397_));
  NAND2_X1  g211(.A1(new_n397_), .A2(G122), .ZN(new_n398_));
  AOI21_X1  g212(.A(new_n211_), .B1(new_n398_), .B2(KEYINPUT37), .ZN(new_n399_));
  INV_X1    g213(.A(G122), .ZN(new_n400_));
  NAND2_X1  g214(.A1(new_n400_), .A2(G116), .ZN(new_n401_));
  NAND2_X1  g215(.A1(new_n401_), .A2(new_n398_), .ZN(new_n402_));
  XNOR2_X1  g216(.A(new_n399_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g217(.A(KEYINPUT34), .ZN(new_n404_));
  NAND3_X1  g218(.A1(new_n404_), .A2(new_n241_), .A3(G128), .ZN(new_n405_));
  AOI21_X1  g219(.A(KEYINPUT34), .B1(new_n238_), .B2(G143), .ZN(new_n406_));
  NOR2_X1   g220(.A1(new_n238_), .A2(G143), .ZN(new_n407_));
  OAI211_X1 g221(.A(new_n190_), .B(new_n405_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g222(.A1(new_n238_), .A2(G143), .ZN(new_n409_));
  NAND2_X1  g223(.A1(new_n409_), .A2(new_n404_), .ZN(new_n410_));
  NAND2_X1  g224(.A1(new_n241_), .A2(G128), .ZN(new_n411_));
  NAND2_X1  g225(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g226(.A1(new_n412_), .A2(new_n405_), .ZN(new_n413_));
  NAND2_X1  g227(.A1(new_n413_), .A2(G134), .ZN(new_n414_));
  AOI21_X1  g228(.A(new_n403_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g229(.A(new_n190_), .B1(new_n411_), .B2(new_n409_), .ZN(new_n416_));
  XNOR2_X1  g230(.A(G116), .B(G122), .ZN(new_n417_));
  NAND2_X1  g231(.A1(new_n417_), .A2(new_n211_), .ZN(new_n418_));
  NOR2_X1   g232(.A1(new_n397_), .A2(G122), .ZN(new_n419_));
  NOR2_X1   g233(.A1(new_n400_), .A2(G116), .ZN(new_n420_));
  OAI21_X1  g234(.A(G107), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g235(.A(new_n416_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g236(.A1(new_n412_), .A2(KEYINPUT35), .A3(new_n190_), .A4(new_n405_), .ZN(new_n423_));
  INV_X1    g237(.A(KEYINPUT35), .ZN(new_n424_));
  NAND2_X1  g238(.A1(new_n408_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g239(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g240(.A(KEYINPUT36), .ZN(new_n427_));
  NAND2_X1  g241(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g242(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT36), .A4(new_n425_), .ZN(new_n429_));
  AOI21_X1  g243(.A(new_n415_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g244(.A1(new_n277_), .A2(G217), .A3(G234), .ZN(new_n431_));
  XNOR2_X1  g245(.A(new_n431_), .B(KEYINPUT33), .ZN(new_n432_));
  NOR2_X1   g246(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g247(.A1(new_n428_), .A2(new_n429_), .ZN(new_n434_));
  INV_X1    g248(.A(new_n415_), .ZN(new_n435_));
  AND3_X1   g249(.A1(new_n434_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  OAI211_X1 g250(.A(new_n395_), .B(new_n396_), .C1(new_n433_), .C2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g251(.A1(new_n437_), .A2(KEYINPUT38), .ZN(new_n438_));
  OAI21_X1  g252(.A(new_n396_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n439_));
  NAND2_X1  g253(.A1(new_n439_), .A2(G478), .ZN(new_n440_));
  XNOR2_X1  g254(.A(new_n438_), .B(new_n440_), .ZN(new_n441_));
  NOR3_X1   g255(.A1(new_n386_), .A2(new_n394_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n443_));
  INV_X1    g257(.A(G113), .ZN(new_n444_));
  INV_X1    g258(.A(G119), .ZN(new_n445_));
  NAND2_X1  g259(.A1(new_n445_), .A2(G116), .ZN(new_n446_));
  NAND2_X1  g260(.A1(new_n397_), .A2(G119), .ZN(new_n447_));
  AOI21_X1  g261(.A(new_n444_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OR2_X1    g262(.A1(new_n448_), .A2(KEYINPUT8), .ZN(new_n449_));
  NOR2_X1   g263(.A1(new_n445_), .A2(G116), .ZN(new_n450_));
  OAI21_X1  g264(.A(new_n446_), .B1(new_n450_), .B2(KEYINPUT4), .ZN(new_n451_));
  OR3_X1    g265(.A1(new_n397_), .A2(KEYINPUT4), .A3(G119), .ZN(new_n452_));
  NAND3_X1  g266(.A1(new_n451_), .A2(new_n444_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g267(.A1(new_n448_), .A2(KEYINPUT8), .ZN(new_n454_));
  NAND3_X1  g268(.A1(new_n449_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g269(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g270(.A(new_n443_), .B1(new_n237_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g271(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n458_));
  NAND3_X1  g272(.A1(new_n458_), .A2(KEYINPUT19), .A3(new_n455_), .ZN(new_n459_));
  OAI211_X1 g273(.A(new_n256_), .B(new_n456_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n460_));
  INV_X1    g274(.A(KEYINPUT20), .ZN(new_n461_));
  NAND2_X1  g275(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g276(.A1(new_n265_), .A2(KEYINPUT20), .A3(new_n256_), .A4(new_n456_), .ZN(new_n463_));
  NAND4_X1  g277(.A1(new_n457_), .A2(new_n459_), .A3(new_n462_), .A4(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465_));
  XOR2_X1   g279(.A(new_n465_), .B(KEYINPUT3), .Z(new_n466_));
  XNOR2_X1  g280(.A(new_n466_), .B(KEYINPUT18), .ZN(new_n467_));
  NAND2_X1  g281(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g282(.A(new_n460_), .ZN(new_n469_));
  INV_X1    g283(.A(KEYINPUT5), .ZN(new_n470_));
  NAND2_X1  g284(.A1(new_n453_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g285(.A1(new_n451_), .A2(KEYINPUT5), .A3(new_n444_), .A4(new_n452_), .ZN(new_n472_));
  NAND2_X1  g286(.A1(new_n451_), .A2(new_n452_), .ZN(new_n473_));
  NAND2_X1  g287(.A1(new_n473_), .A2(G113), .ZN(new_n474_));
  NAND3_X1  g288(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  AOI22_X1  g289(.A1(new_n469_), .A2(KEYINPUT13), .B1(new_n475_), .B2(new_n268_), .ZN(new_n476_));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477_));
  INV_X1    g291(.A(new_n466_), .ZN(new_n478_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n479_));
  NAND2_X1  g293(.A1(new_n460_), .A2(new_n479_), .ZN(new_n480_));
  NAND4_X1  g294(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  NAND4_X1  g295(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n256_), .A4(new_n456_), .ZN(new_n482_));
  NAND2_X1  g296(.A1(new_n268_), .A2(new_n475_), .ZN(new_n483_));
  NAND4_X1  g297(.A1(new_n480_), .A2(new_n482_), .A3(new_n478_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g298(.A1(new_n484_), .A2(KEYINPUT17), .ZN(new_n485_));
  MUX2_X1   g299(.A(new_n254_), .B(new_n271_), .S(G125), .Z(new_n486_));
  AND2_X1   g300(.A1(new_n277_), .A2(G224), .ZN(new_n487_));
  NOR2_X1   g301(.A1(new_n487_), .A2(KEYINPUT16), .ZN(new_n488_));
  XNOR2_X1  g302(.A(new_n486_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g303(.A(new_n489_), .ZN(new_n490_));
  NAND4_X1  g304(.A1(new_n468_), .A2(new_n481_), .A3(new_n485_), .A4(new_n490_), .ZN(new_n491_));
  NAND2_X1  g305(.A1(new_n491_), .A2(KEYINPUT21), .ZN(new_n492_));
  AOI21_X1  g306(.A(new_n489_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n493_));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n494_));
  NAND4_X1  g308(.A1(new_n493_), .A2(new_n494_), .A3(new_n481_), .A4(new_n485_), .ZN(new_n495_));
  AND2_X1   g309(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497_));
  XNOR2_X1  g311(.A(new_n497_), .B(KEYINPUT22), .ZN(new_n498_));
  NAND4_X1  g312(.A1(new_n476_), .A2(KEYINPUT14), .A3(new_n478_), .A4(new_n480_), .ZN(new_n499_));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n500_));
  NAND2_X1  g314(.A1(new_n484_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g315(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g316(.A1(new_n480_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n503_));
  AOI21_X1  g317(.A(KEYINPUT15), .B1(new_n503_), .B2(new_n466_), .ZN(new_n504_));
  NAND3_X1  g318(.A1(new_n503_), .A2(KEYINPUT15), .A3(new_n466_), .ZN(new_n505_));
  INV_X1    g319(.A(new_n505_), .ZN(new_n506_));
  OAI21_X1  g320(.A(new_n502_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g321(.A(new_n486_), .B(new_n487_), .ZN(new_n508_));
  INV_X1    g322(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g323(.A(new_n188_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g324(.A1(new_n496_), .A2(KEYINPUT23), .A3(new_n498_), .A4(new_n510_), .ZN(new_n511_));
  NAND2_X1  g325(.A1(new_n498_), .A2(KEYINPUT23), .ZN(new_n512_));
  OR2_X1    g326(.A1(new_n498_), .A2(KEYINPUT23), .ZN(new_n513_));
  NAND2_X1  g327(.A1(new_n492_), .A2(new_n495_), .ZN(new_n514_));
  NAND2_X1  g328(.A1(new_n503_), .A2(new_n466_), .ZN(new_n515_));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n516_));
  NAND2_X1  g330(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g331(.A1(new_n517_), .A2(new_n505_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n518_));
  OAI21_X1  g332(.A(new_n396_), .B1(new_n518_), .B2(new_n508_), .ZN(new_n519_));
  OAI211_X1 g333(.A(new_n512_), .B(new_n513_), .C1(new_n514_), .C2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g334(.A(G214), .B1(G237), .B2(G902), .ZN(new_n521_));
  NAND3_X1  g335(.A1(new_n511_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g336(.A1(new_n522_), .A2(KEYINPUT24), .ZN(new_n523_));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n524_));
  NAND4_X1  g338(.A1(new_n511_), .A2(new_n520_), .A3(new_n524_), .A4(new_n521_), .ZN(new_n525_));
  NAND2_X1  g339(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  AND3_X1   g340(.A1(new_n320_), .A2(new_n442_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n528_));
  INV_X1    g342(.A(G472), .ZN(new_n529_));
  NAND2_X1  g343(.A1(new_n206_), .A2(new_n271_), .ZN(new_n530_));
  NAND2_X1  g344(.A1(new_n530_), .A2(KEYINPUT60), .ZN(new_n531_));
  INV_X1    g345(.A(KEYINPUT60), .ZN(new_n532_));
  NAND3_X1  g346(.A1(new_n206_), .A2(new_n532_), .A3(new_n271_), .ZN(new_n533_));
  NAND2_X1  g347(.A1(new_n195_), .A2(KEYINPUT59), .ZN(new_n534_));
  NAND2_X1  g348(.A1(new_n191_), .A2(KEYINPUT58), .ZN(new_n535_));
  NAND2_X1  g349(.A1(new_n535_), .A2(new_n197_), .ZN(new_n536_));
  NOR2_X1   g350(.A1(new_n191_), .A2(KEYINPUT58), .ZN(new_n537_));
  OAI21_X1  g351(.A(G131), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g352(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g353(.A(KEYINPUT59), .ZN(new_n540_));
  OAI211_X1 g354(.A(new_n254_), .B(new_n539_), .C1(new_n540_), .C2(new_n538_), .ZN(new_n541_));
  NAND3_X1  g355(.A1(new_n531_), .A2(new_n533_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g356(.A1(new_n542_), .A2(KEYINPUT63), .ZN(new_n543_));
  INV_X1    g357(.A(KEYINPUT57), .ZN(new_n544_));
  XNOR2_X1  g358(.A(new_n475_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g359(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g360(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g361(.A1(new_n324_), .A2(G210), .ZN(new_n548_));
  XNOR2_X1  g362(.A(KEYINPUT56), .B(G101), .ZN(new_n549_));
  XNOR2_X1  g363(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g364(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g365(.A1(new_n542_), .A2(KEYINPUT63), .A3(new_n545_), .ZN(new_n552_));
  NAND3_X1  g366(.A1(new_n547_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g367(.A1(new_n542_), .A2(new_n545_), .ZN(new_n554_));
  NAND2_X1  g368(.A1(new_n554_), .A2(KEYINPUT61), .ZN(new_n555_));
  INV_X1    g369(.A(new_n542_), .ZN(new_n556_));
  NAND2_X1  g370(.A1(new_n556_), .A2(new_n546_), .ZN(new_n557_));
  INV_X1    g371(.A(KEYINPUT61), .ZN(new_n558_));
  NAND3_X1  g372(.A1(new_n542_), .A2(new_n558_), .A3(new_n545_), .ZN(new_n559_));
  NAND3_X1  g373(.A1(new_n555_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  AOI22_X1  g374(.A1(KEYINPUT65), .A2(new_n553_), .B1(new_n560_), .B2(new_n550_), .ZN(new_n561_));
  AND3_X1   g375(.A1(new_n560_), .A2(KEYINPUT65), .A3(new_n550_), .ZN(new_n562_));
  OAI211_X1 g376(.A(new_n529_), .B(new_n396_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g377(.A(KEYINPUT66), .ZN(new_n564_));
  NAND2_X1  g378(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g379(.A1(new_n560_), .A2(new_n550_), .ZN(new_n566_));
  NAND2_X1  g380(.A1(new_n553_), .A2(KEYINPUT65), .ZN(new_n567_));
  NAND2_X1  g381(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g382(.A1(new_n560_), .A2(KEYINPUT65), .A3(new_n550_), .ZN(new_n569_));
  NAND2_X1  g383(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g384(.A1(new_n570_), .A2(KEYINPUT66), .A3(new_n529_), .A4(new_n396_), .ZN(new_n571_));
  NOR2_X1   g385(.A1(new_n396_), .A2(new_n529_), .ZN(new_n572_));
  INV_X1    g386(.A(new_n572_), .ZN(new_n573_));
  NAND4_X1  g387(.A1(new_n555_), .A2(new_n557_), .A3(new_n559_), .A4(new_n551_), .ZN(new_n574_));
  INV_X1    g388(.A(KEYINPUT62), .ZN(new_n575_));
  NAND2_X1  g389(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g390(.A1(new_n576_), .A2(G472), .ZN(new_n577_));
  INV_X1    g391(.A(new_n552_), .ZN(new_n578_));
  AOI21_X1  g392(.A(new_n545_), .B1(new_n542_), .B2(KEYINPUT63), .ZN(new_n579_));
  OAI21_X1  g393(.A(new_n550_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g394(.A(new_n575_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n581_));
  OAI21_X1  g395(.A(new_n573_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g396(.A(KEYINPUT64), .ZN(new_n583_));
  NAND2_X1  g397(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g398(.A(KEYINPUT64), .B(new_n573_), .C1(new_n577_), .C2(new_n581_), .ZN(new_n585_));
  AOI22_X1  g399(.A1(new_n565_), .A2(new_n571_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g400(.A(KEYINPUT55), .ZN(new_n587_));
  XNOR2_X1  g401(.A(KEYINPUT53), .B(G110), .ZN(new_n588_));
  INV_X1    g402(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g403(.A(G119), .B(G128), .ZN(new_n590_));
  NAND2_X1  g404(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g405(.A(G110), .ZN(new_n592_));
  OAI211_X1 g406(.A(new_n346_), .B(new_n591_), .C1(new_n592_), .C2(new_n590_), .ZN(new_n593_));
  XOR2_X1   g407(.A(new_n344_), .B(KEYINPUT52), .Z(new_n594_));
  NAND2_X1  g408(.A1(new_n590_), .A2(G110), .ZN(new_n595_));
  OAI211_X1 g409(.A(new_n345_), .B(new_n595_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n596_));
  OAI21_X1  g410(.A(new_n593_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g411(.A1(new_n281_), .A2(G221), .A3(G234), .ZN(new_n598_));
  XNOR2_X1  g412(.A(new_n598_), .B(new_n192_), .ZN(new_n599_));
  NAND2_X1  g413(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g414(.A1(new_n600_), .A2(KEYINPUT54), .ZN(new_n601_));
  OR2_X1    g415(.A1(new_n597_), .A2(new_n599_), .ZN(new_n602_));
  XNOR2_X1  g416(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g417(.A(new_n603_), .ZN(new_n604_));
  OAI21_X1  g418(.A(new_n587_), .B1(new_n604_), .B2(new_n188_), .ZN(new_n605_));
  INV_X1    g419(.A(G217), .ZN(new_n606_));
  AOI21_X1  g420(.A(new_n606_), .B1(new_n396_), .B2(G234), .ZN(new_n607_));
  NAND3_X1  g421(.A1(new_n603_), .A2(KEYINPUT55), .A3(new_n396_), .ZN(new_n608_));
  NAND3_X1  g422(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g423(.A(new_n607_), .ZN(new_n610_));
  NAND3_X1  g424(.A1(new_n603_), .A2(new_n396_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g425(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g426(.A(new_n528_), .B1(new_n586_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g427(.A1(new_n565_), .A2(new_n571_), .ZN(new_n614_));
  NAND2_X1  g428(.A1(new_n584_), .A2(new_n585_), .ZN(new_n615_));
  NAND2_X1  g429(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g430(.A(new_n612_), .ZN(new_n617_));
  NAND3_X1  g431(.A1(new_n616_), .A2(KEYINPUT67), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g432(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g433(.A1(new_n527_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g434(.A(new_n620_), .B(G101), .ZN(G3));
  AND2_X1   g435(.A1(new_n526_), .A2(new_n392_), .ZN(new_n622_));
  INV_X1    g436(.A(new_n437_), .ZN(new_n623_));
  INV_X1    g437(.A(KEYINPUT69), .ZN(new_n624_));
  XOR2_X1   g438(.A(new_n432_), .B(KEYINPUT68), .Z(new_n625_));
  INV_X1    g439(.A(new_n625_), .ZN(new_n626_));
  NOR3_X1   g440(.A1(new_n430_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g441(.A1(new_n430_), .A2(new_n432_), .ZN(new_n628_));
  NAND2_X1  g442(.A1(new_n628_), .A2(KEYINPUT69), .ZN(new_n629_));
  NAND2_X1  g443(.A1(new_n434_), .A2(new_n435_), .ZN(new_n630_));
  NAND2_X1  g444(.A1(new_n630_), .A2(new_n625_), .ZN(new_n631_));
  AOI21_X1  g445(.A(new_n627_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g446(.A(G478), .B1(new_n632_), .B2(new_n188_), .ZN(new_n633_));
  AOI21_X1  g447(.A(new_n623_), .B1(new_n633_), .B2(KEYINPUT70), .ZN(new_n634_));
  INV_X1    g448(.A(KEYINPUT70), .ZN(new_n635_));
  OAI211_X1 g449(.A(new_n635_), .B(G478), .C1(new_n632_), .C2(new_n188_), .ZN(new_n636_));
  AOI21_X1  g450(.A(KEYINPUT71), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g451(.A(new_n631_), .B1(new_n436_), .B2(new_n624_), .ZN(new_n638_));
  INV_X1    g452(.A(new_n627_), .ZN(new_n639_));
  AOI21_X1  g453(.A(new_n188_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g454(.A(KEYINPUT70), .B1(new_n640_), .B2(new_n395_), .ZN(new_n641_));
  AND4_X1   g455(.A1(KEYINPUT71), .A2(new_n641_), .A3(new_n437_), .A4(new_n636_), .ZN(new_n642_));
  NOR2_X1   g456(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g457(.A1(new_n385_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g458(.A1(new_n622_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g459(.A(new_n188_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n646_));
  INV_X1    g460(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g461(.A1(new_n647_), .A2(KEYINPUT72), .A3(G472), .ZN(new_n648_));
  INV_X1    g462(.A(KEYINPUT72), .ZN(new_n649_));
  OAI21_X1  g463(.A(new_n649_), .B1(new_n646_), .B2(new_n529_), .ZN(new_n650_));
  NAND2_X1  g464(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g465(.A1(new_n570_), .A2(new_n529_), .A3(new_n372_), .ZN(new_n652_));
  INV_X1    g466(.A(KEYINPUT73), .ZN(new_n653_));
  NAND2_X1  g467(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g468(.A1(new_n570_), .A2(KEYINPUT73), .A3(new_n529_), .A4(new_n372_), .ZN(new_n655_));
  NAND2_X1  g469(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g470(.A1(new_n651_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g471(.A1(new_n657_), .A2(new_n612_), .ZN(new_n658_));
  AND2_X1   g472(.A1(new_n320_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g473(.A1(new_n645_), .A2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g474(.A(new_n660_), .B(G104), .ZN(G6));
  AND2_X1   g475(.A1(new_n362_), .A2(new_n365_), .ZN(new_n662_));
  INV_X1    g476(.A(new_n367_), .ZN(new_n663_));
  OAI21_X1  g477(.A(new_n396_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI22_X1  g478(.A1(new_n664_), .A2(G475), .B1(new_n383_), .B2(new_n384_), .ZN(new_n665_));
  NAND2_X1  g479(.A1(new_n665_), .A2(new_n441_), .ZN(new_n666_));
  INV_X1    g480(.A(new_n666_), .ZN(new_n667_));
  AND2_X1   g481(.A1(new_n622_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g482(.A1(new_n668_), .A2(new_n659_), .ZN(new_n669_));
  XNOR2_X1  g483(.A(new_n669_), .B(G107), .ZN(G9));
  INV_X1    g484(.A(KEYINPUT74), .ZN(new_n671_));
  NAND2_X1  g485(.A1(new_n602_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g486(.A(new_n672_), .B(new_n600_), .ZN(new_n673_));
  NAND2_X1  g487(.A1(new_n673_), .A2(new_n610_), .ZN(new_n674_));
  AOI21_X1  g488(.A(new_n188_), .B1(new_n674_), .B2(KEYINPUT75), .ZN(new_n675_));
  OAI21_X1  g489(.A(new_n675_), .B1(KEYINPUT75), .B2(new_n674_), .ZN(new_n676_));
  NAND2_X1  g490(.A1(new_n676_), .A2(new_n609_), .ZN(new_n677_));
  AND3_X1   g491(.A1(new_n651_), .A2(new_n656_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g492(.A1(new_n527_), .A2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g493(.A(KEYINPUT76), .B(G110), .Z(new_n680_));
  XNOR2_X1  g494(.A(new_n679_), .B(new_n680_), .ZN(G12));
  XOR2_X1   g495(.A(KEYINPUT77), .B(G900), .Z(new_n682_));
  NAND3_X1  g496(.A1(new_n682_), .A2(G953), .A3(new_n389_), .ZN(new_n683_));
  XOR2_X1   g497(.A(new_n683_), .B(KEYINPUT78), .Z(new_n684_));
  NOR2_X1   g498(.A1(new_n684_), .A2(new_n388_), .ZN(new_n685_));
  NOR2_X1   g499(.A1(new_n666_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g500(.A1(new_n526_), .A2(new_n686_), .ZN(new_n687_));
  AOI22_X1  g501(.A1(new_n614_), .A2(new_n615_), .B1(new_n609_), .B2(new_n676_), .ZN(new_n688_));
  AOI21_X1  g502(.A(new_n318_), .B1(new_n317_), .B2(new_n307_), .ZN(new_n689_));
  AOI211_X1 g503(.A(KEYINPUT32), .B(new_n308_), .C1(new_n311_), .C2(new_n316_), .ZN(new_n690_));
  OAI21_X1  g504(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g505(.A(KEYINPUT79), .B1(new_n687_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g506(.A(new_n686_), .ZN(new_n693_));
  AOI21_X1  g507(.A(new_n693_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n694_));
  NAND2_X1  g508(.A1(new_n616_), .A2(new_n677_), .ZN(new_n695_));
  AOI21_X1  g509(.A(new_n695_), .B1(new_n309_), .B2(new_n319_), .ZN(new_n696_));
  INV_X1    g510(.A(KEYINPUT79), .ZN(new_n697_));
  NAND3_X1  g511(.A1(new_n694_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g512(.A1(new_n692_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g513(.A(KEYINPUT80), .B(G128), .ZN(new_n700_));
  XNOR2_X1  g514(.A(new_n699_), .B(new_n700_), .ZN(G30));
  INV_X1    g515(.A(new_n553_), .ZN(new_n702_));
  XOR2_X1   g516(.A(new_n557_), .B(KEYINPUT81), .Z(new_n703_));
  NAND3_X1  g517(.A1(new_n703_), .A2(new_n559_), .A3(new_n555_), .ZN(new_n704_));
  AOI21_X1  g518(.A(new_n702_), .B1(new_n704_), .B2(new_n550_), .ZN(new_n705_));
  OAI21_X1  g519(.A(G472), .B1(new_n705_), .B2(G902), .ZN(new_n706_));
  AND2_X1   g520(.A1(new_n706_), .A2(new_n614_), .ZN(new_n707_));
  NOR2_X1   g521(.A1(new_n707_), .A2(new_n677_), .ZN(new_n708_));
  INV_X1    g522(.A(new_n441_), .ZN(new_n709_));
  NOR2_X1   g523(.A1(new_n385_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g524(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g525(.A(new_n685_), .ZN(new_n712_));
  NAND3_X1  g526(.A1(new_n317_), .A2(new_n307_), .A3(new_n712_), .ZN(new_n713_));
  AND2_X1   g527(.A1(new_n713_), .A2(KEYINPUT82), .ZN(new_n714_));
  NOR2_X1   g528(.A1(new_n713_), .A2(KEYINPUT82), .ZN(new_n715_));
  NOR4_X1   g529(.A1(new_n711_), .A2(new_n714_), .A3(new_n715_), .A4(new_n522_), .ZN(new_n716_));
  XNOR2_X1  g530(.A(new_n716_), .B(new_n241_), .ZN(G45));
  NAND2_X1  g531(.A1(new_n373_), .A2(KEYINPUT48), .ZN(new_n718_));
  NAND3_X1  g532(.A1(new_n718_), .A2(G475), .A3(new_n376_), .ZN(new_n719_));
  NAND2_X1  g533(.A1(new_n383_), .A2(new_n384_), .ZN(new_n720_));
  AOI211_X1 g534(.A(new_n685_), .B(new_n643_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g535(.A1(new_n320_), .A2(new_n526_), .A3(new_n688_), .A4(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g536(.A(new_n722_), .B(G146), .ZN(G48));
  INV_X1    g537(.A(new_n619_), .ZN(new_n724_));
  AOI21_X1  g538(.A(G469), .B1(new_n312_), .B2(new_n372_), .ZN(new_n725_));
  NOR2_X1   g539(.A1(new_n188_), .A2(new_n187_), .ZN(new_n726_));
  AOI21_X1  g540(.A(new_n725_), .B1(new_n303_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g541(.A(KEYINPUT83), .B1(new_n727_), .B2(new_n308_), .ZN(new_n728_));
  INV_X1    g542(.A(KEYINPUT83), .ZN(new_n729_));
  AND3_X1   g543(.A1(new_n314_), .A2(new_n315_), .A3(new_n726_), .ZN(new_n730_));
  OAI211_X1 g544(.A(new_n729_), .B(new_n307_), .C1(new_n730_), .C2(new_n725_), .ZN(new_n731_));
  NAND2_X1  g545(.A1(new_n728_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g546(.A(new_n732_), .ZN(new_n733_));
  NOR2_X1   g547(.A1(new_n724_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g548(.A1(new_n645_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g549(.A(new_n735_), .B(G113), .ZN(G15));
  NAND2_X1  g550(.A1(new_n668_), .A2(new_n734_), .ZN(new_n737_));
  NAND2_X1  g551(.A1(new_n737_), .A2(KEYINPUT84), .ZN(new_n738_));
  INV_X1    g552(.A(KEYINPUT84), .ZN(new_n739_));
  NAND3_X1  g553(.A1(new_n668_), .A2(new_n739_), .A3(new_n734_), .ZN(new_n740_));
  NAND2_X1  g554(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g555(.A(new_n741_), .B(G116), .ZN(G18));
  NAND4_X1  g556(.A1(new_n442_), .A2(new_n526_), .A3(new_n688_), .A4(new_n732_), .ZN(new_n743_));
  XOR2_X1   g557(.A(KEYINPUT85), .B(G119), .Z(new_n744_));
  XNOR2_X1  g558(.A(new_n743_), .B(new_n744_), .ZN(G21));
  NOR2_X1   g559(.A1(new_n522_), .A2(new_n394_), .ZN(new_n746_));
  XNOR2_X1  g560(.A(new_n746_), .B(KEYINPUT86), .ZN(new_n747_));
  NAND4_X1  g561(.A1(new_n747_), .A2(new_n658_), .A3(new_n710_), .A4(new_n732_), .ZN(new_n748_));
  XNOR2_X1  g562(.A(new_n748_), .B(G122), .ZN(G24));
  NAND4_X1  g563(.A1(new_n732_), .A2(new_n526_), .A3(new_n678_), .A4(new_n721_), .ZN(new_n750_));
  XOR2_X1   g564(.A(KEYINPUT87), .B(G125), .Z(new_n751_));
  XNOR2_X1  g565(.A(new_n750_), .B(new_n751_), .ZN(G27));
  NAND2_X1  g566(.A1(new_n511_), .A2(new_n520_), .ZN(new_n753_));
  NAND2_X1  g567(.A1(new_n753_), .A2(new_n521_), .ZN(new_n754_));
  INV_X1    g568(.A(new_n754_), .ZN(new_n755_));
  NAND2_X1  g569(.A1(new_n320_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g570(.A1(new_n724_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g571(.A1(new_n757_), .A2(new_n721_), .ZN(new_n758_));
  XNOR2_X1  g572(.A(new_n758_), .B(G131), .ZN(G33));
  NAND2_X1  g573(.A1(new_n757_), .A2(new_n686_), .ZN(new_n760_));
  XNOR2_X1  g574(.A(new_n760_), .B(G134), .ZN(G36));
  INV_X1    g575(.A(new_n643_), .ZN(new_n762_));
  AND2_X1   g576(.A1(new_n762_), .A2(new_n665_), .ZN(new_n763_));
  AND2_X1   g577(.A1(new_n763_), .A2(new_n677_), .ZN(new_n764_));
  AND3_X1   g578(.A1(new_n314_), .A2(new_n315_), .A3(new_n304_), .ZN(new_n765_));
  NAND2_X1  g579(.A1(new_n261_), .A2(new_n273_), .ZN(new_n766_));
  INV_X1    g580(.A(KEYINPUT88), .ZN(new_n767_));
  AOI21_X1  g581(.A(new_n284_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g582(.A(new_n768_), .B1(new_n767_), .B2(new_n766_), .ZN(new_n769_));
  NAND3_X1  g583(.A1(new_n293_), .A2(KEYINPUT89), .A3(new_n284_), .ZN(new_n770_));
  OAI21_X1  g584(.A(new_n770_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n771_));
  AOI21_X1  g585(.A(KEYINPUT89), .B1(new_n293_), .B2(new_n284_), .ZN(new_n772_));
  OAI21_X1  g586(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g587(.A(new_n187_), .B1(new_n773_), .B2(new_n372_), .ZN(new_n774_));
  OAI211_X1 g588(.A(new_n307_), .B(new_n712_), .C1(new_n765_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g589(.A(new_n775_), .ZN(new_n776_));
  NAND4_X1  g590(.A1(new_n764_), .A2(new_n657_), .A3(new_n755_), .A4(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g591(.A(new_n777_), .B(G137), .ZN(G39));
  NOR2_X1   g592(.A1(new_n765_), .A2(new_n774_), .ZN(new_n779_));
  OR3_X1    g593(.A1(new_n779_), .A2(KEYINPUT90), .A3(new_n308_), .ZN(new_n780_));
  OAI21_X1  g594(.A(KEYINPUT90), .B1(new_n779_), .B2(new_n308_), .ZN(new_n781_));
  NAND2_X1  g595(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR3_X1   g596(.A1(new_n754_), .A2(new_n617_), .A3(new_n616_), .ZN(new_n783_));
  NAND3_X1  g597(.A1(new_n782_), .A2(new_n721_), .A3(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g598(.A(new_n784_), .B(G140), .ZN(G42));
  NAND3_X1  g599(.A1(new_n707_), .A2(new_n753_), .A3(new_n385_), .ZN(new_n786_));
  XNOR2_X1  g600(.A(new_n786_), .B(KEYINPUT95), .ZN(new_n787_));
  NAND3_X1  g601(.A1(new_n762_), .A2(new_n617_), .A3(new_n521_), .ZN(new_n788_));
  NOR4_X1   g602(.A1(new_n787_), .A2(new_n308_), .A3(new_n727_), .A4(new_n788_), .ZN(new_n789_));
  NOR3_X1   g603(.A1(new_n789_), .A2(G952), .A3(G953), .ZN(new_n790_));
  NAND2_X1  g604(.A1(new_n763_), .A2(new_n388_), .ZN(new_n791_));
  XNOR2_X1  g605(.A(new_n791_), .B(KEYINPUT93), .ZN(new_n792_));
  NOR3_X1   g606(.A1(new_n792_), .A2(new_n612_), .A3(new_n657_), .ZN(new_n793_));
  XNOR2_X1  g607(.A(new_n793_), .B(KEYINPUT96), .ZN(new_n794_));
  NAND3_X1  g608(.A1(new_n794_), .A2(new_n526_), .A3(new_n732_), .ZN(new_n795_));
  XOR2_X1   g609(.A(new_n795_), .B(KEYINPUT97), .Z(new_n796_));
  INV_X1    g610(.A(new_n782_), .ZN(new_n797_));
  OAI21_X1  g611(.A(new_n308_), .B1(new_n730_), .B2(new_n725_), .ZN(new_n798_));
  AOI21_X1  g612(.A(new_n754_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g613(.A(new_n521_), .B1(new_n511_), .B2(new_n520_), .ZN(new_n800_));
  XNOR2_X1  g614(.A(new_n800_), .B(KEYINPUT98), .ZN(new_n801_));
  NOR2_X1   g615(.A1(new_n733_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g616(.A(new_n794_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g617(.A1(new_n755_), .A2(new_n617_), .A3(new_n388_), .A4(new_n707_), .ZN(new_n804_));
  NOR4_X1   g618(.A1(new_n804_), .A2(new_n733_), .A3(new_n386_), .A4(new_n762_), .ZN(new_n805_));
  INV_X1    g619(.A(KEYINPUT99), .ZN(new_n806_));
  NOR2_X1   g620(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR3_X1   g621(.A1(new_n792_), .A2(new_n733_), .A3(new_n754_), .ZN(new_n808_));
  AOI211_X1 g622(.A(new_n789_), .B(new_n807_), .C1(new_n678_), .C2(new_n808_), .ZN(new_n809_));
  AND2_X1   g623(.A1(new_n808_), .A2(new_n619_), .ZN(new_n810_));
  NAND2_X1  g624(.A1(new_n810_), .A2(KEYINPUT94), .ZN(new_n811_));
  NAND2_X1  g625(.A1(new_n281_), .A2(G952), .ZN(new_n812_));
  AOI21_X1  g626(.A(new_n812_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n813_));
  NAND4_X1  g627(.A1(new_n803_), .A2(new_n809_), .A3(new_n811_), .A4(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g628(.A(new_n644_), .B(KEYINPUT91), .ZN(new_n815_));
  NOR3_X1   g629(.A1(new_n815_), .A2(new_n733_), .A3(new_n804_), .ZN(new_n816_));
  XNOR2_X1  g630(.A(new_n816_), .B(KEYINPUT92), .ZN(new_n817_));
  OAI21_X1  g631(.A(new_n817_), .B1(KEYINPUT94), .B2(new_n810_), .ZN(new_n818_));
  NOR3_X1   g632(.A1(new_n796_), .A2(new_n814_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g633(.A1(new_n722_), .A2(new_n750_), .ZN(new_n820_));
  XNOR2_X1  g634(.A(new_n820_), .B(KEYINPUT104), .ZN(new_n821_));
  AOI21_X1  g635(.A(new_n711_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n822_));
  AOI21_X1  g636(.A(new_n685_), .B1(new_n309_), .B2(new_n319_), .ZN(new_n823_));
  AOI22_X1  g637(.A1(new_n822_), .A2(new_n823_), .B1(new_n692_), .B2(new_n698_), .ZN(new_n824_));
  NAND2_X1  g638(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  OR2_X1    g639(.A1(new_n825_), .A2(KEYINPUT105), .ZN(new_n826_));
  NAND2_X1  g640(.A1(new_n825_), .A2(KEYINPUT105), .ZN(new_n827_));
  NAND2_X1  g641(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OR2_X1    g642(.A1(new_n756_), .A2(KEYINPUT100), .ZN(new_n829_));
  NAND2_X1  g643(.A1(new_n756_), .A2(KEYINPUT100), .ZN(new_n830_));
  NAND4_X1  g644(.A1(new_n829_), .A2(new_n678_), .A3(new_n721_), .A4(new_n830_), .ZN(new_n831_));
  NOR2_X1   g645(.A1(new_n386_), .A2(new_n441_), .ZN(new_n832_));
  AOI211_X1 g646(.A(new_n754_), .B(new_n695_), .C1(new_n832_), .C2(KEYINPUT101), .ZN(new_n833_));
  OAI211_X1 g647(.A(new_n833_), .B(new_n823_), .C1(KEYINPUT101), .C2(new_n832_), .ZN(new_n834_));
  AOI21_X1  g648(.A(new_n754_), .B1(new_n309_), .B2(new_n319_), .ZN(new_n835_));
  OAI211_X1 g649(.A(new_n835_), .B(new_n619_), .C1(new_n686_), .C2(new_n721_), .ZN(new_n836_));
  OR2_X1    g650(.A1(new_n836_), .A2(KEYINPUT102), .ZN(new_n837_));
  NAND3_X1  g651(.A1(new_n831_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g652(.A1(new_n836_), .A2(KEYINPUT102), .ZN(new_n839_));
  INV_X1    g653(.A(new_n839_), .ZN(new_n840_));
  OR3_X1    g654(.A1(new_n838_), .A2(KEYINPUT103), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g655(.A(KEYINPUT103), .B1(new_n838_), .B2(new_n840_), .ZN(new_n842_));
  NAND2_X1  g656(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AND4_X1   g657(.A1(new_n620_), .A2(new_n660_), .A3(new_n669_), .A4(new_n679_), .ZN(new_n844_));
  AND3_X1   g658(.A1(new_n735_), .A2(new_n743_), .A3(new_n748_), .ZN(new_n845_));
  NAND3_X1  g659(.A1(new_n844_), .A2(new_n741_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g660(.A(new_n846_), .ZN(new_n847_));
  NAND3_X1  g661(.A1(new_n828_), .A2(new_n843_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g662(.A1(new_n848_), .A2(KEYINPUT106), .ZN(new_n849_));
  AOI21_X1  g663(.A(new_n846_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n850_));
  INV_X1    g664(.A(KEYINPUT106), .ZN(new_n851_));
  NAND3_X1  g665(.A1(new_n850_), .A2(new_n851_), .A3(new_n843_), .ZN(new_n852_));
  NAND2_X1  g666(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g667(.A(new_n790_), .B1(new_n819_), .B2(new_n853_), .ZN(G75));
  NOR2_X1   g668(.A1(new_n281_), .A2(G952), .ZN(new_n855_));
  INV_X1    g669(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g670(.A(new_n396_), .B1(new_n850_), .B2(new_n843_), .ZN(new_n857_));
  NAND2_X1  g671(.A1(new_n857_), .A2(new_n498_), .ZN(new_n858_));
  XNOR2_X1  g672(.A(new_n507_), .B(KEYINPUT108), .ZN(new_n859_));
  XOR2_X1   g673(.A(new_n508_), .B(KEYINPUT107), .Z(new_n860_));
  XNOR2_X1  g674(.A(new_n859_), .B(new_n860_), .ZN(new_n861_));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862_));
  NAND2_X1  g676(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g677(.A(new_n856_), .B1(new_n858_), .B2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g678(.A(new_n861_), .B(KEYINPUT109), .ZN(new_n865_));
  AOI21_X1  g679(.A(new_n864_), .B1(new_n858_), .B2(new_n865_), .ZN(G51));
  NAND2_X1  g680(.A1(G469), .A2(G902), .ZN(new_n867_));
  OAI21_X1  g681(.A(new_n303_), .B1(new_n853_), .B2(new_n867_), .ZN(new_n868_));
  OR2_X1    g682(.A1(new_n773_), .A2(new_n867_), .ZN(new_n869_));
  INV_X1    g683(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g684(.A1(new_n848_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g685(.A(new_n855_), .B1(new_n868_), .B2(new_n871_), .ZN(G54));
  AOI211_X1 g686(.A(new_n321_), .B(new_n372_), .C1(new_n850_), .C2(new_n843_), .ZN(new_n873_));
  NAND2_X1  g687(.A1(new_n383_), .A2(KEYINPUT110), .ZN(new_n874_));
  INV_X1    g688(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g689(.A(new_n855_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g690(.A(KEYINPUT111), .ZN(new_n877_));
  OAI211_X1 g691(.A(new_n876_), .B(new_n877_), .C1(new_n875_), .C2(new_n873_), .ZN(new_n878_));
  NOR2_X1   g692(.A1(new_n873_), .A2(new_n875_), .ZN(new_n879_));
  NAND3_X1  g693(.A1(new_n848_), .A2(G475), .A3(G902), .ZN(new_n880_));
  OAI21_X1  g694(.A(new_n856_), .B1(new_n880_), .B2(new_n874_), .ZN(new_n881_));
  OAI21_X1  g695(.A(KEYINPUT111), .B1(new_n879_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g696(.A1(new_n878_), .A2(new_n882_), .ZN(G60));
  NOR2_X1   g697(.A1(new_n395_), .A2(new_n372_), .ZN(new_n884_));
  NAND3_X1  g698(.A1(new_n849_), .A2(new_n852_), .A3(new_n884_), .ZN(new_n885_));
  OAI21_X1  g699(.A(new_n856_), .B1(new_n885_), .B2(new_n632_), .ZN(new_n886_));
  AOI21_X1  g700(.A(new_n886_), .B1(new_n632_), .B2(new_n885_), .ZN(G63));
  INV_X1    g701(.A(new_n673_), .ZN(new_n888_));
  NAND4_X1  g702(.A1(new_n848_), .A2(G217), .A3(new_n188_), .A4(new_n888_), .ZN(new_n889_));
  NAND2_X1  g703(.A1(new_n889_), .A2(KEYINPUT112), .ZN(new_n890_));
  INV_X1    g704(.A(KEYINPUT112), .ZN(new_n891_));
  NAND4_X1  g705(.A1(new_n857_), .A2(new_n891_), .A3(G217), .A4(new_n888_), .ZN(new_n892_));
  AND2_X1   g706(.A1(new_n857_), .A2(G217), .ZN(new_n893_));
  OAI211_X1 g707(.A(new_n890_), .B(new_n892_), .C1(new_n893_), .C2(new_n604_), .ZN(new_n894_));
  AND2_X1   g708(.A1(new_n894_), .A2(new_n856_), .ZN(G66));
  NAND2_X1  g709(.A1(new_n846_), .A2(new_n277_), .ZN(new_n896_));
  NAND2_X1  g710(.A1(new_n896_), .A2(KEYINPUT113), .ZN(new_n897_));
  OAI21_X1  g711(.A(new_n859_), .B1(G898), .B2(new_n281_), .ZN(new_n898_));
  INV_X1    g712(.A(new_n898_), .ZN(new_n899_));
  INV_X1    g713(.A(KEYINPUT113), .ZN(new_n900_));
  NAND3_X1  g714(.A1(new_n846_), .A2(new_n900_), .A3(new_n277_), .ZN(new_n901_));
  NAND3_X1  g715(.A1(new_n897_), .A2(new_n899_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n903_));
  AND2_X1   g717(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g718(.A(new_n901_), .ZN(new_n905_));
  AOI21_X1  g719(.A(new_n900_), .B1(new_n846_), .B2(new_n277_), .ZN(new_n906_));
  OAI21_X1  g720(.A(new_n898_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g721(.A(KEYINPUT114), .ZN(new_n908_));
  NOR2_X1   g722(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g723(.A1(new_n902_), .A2(new_n903_), .ZN(new_n910_));
  NOR3_X1   g724(.A1(new_n904_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  AOI21_X1  g725(.A(new_n277_), .B1(G224), .B2(G898), .ZN(new_n912_));
  AOI21_X1  g726(.A(new_n912_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n913_));
  AOI22_X1  g727(.A1(new_n911_), .A2(new_n913_), .B1(new_n912_), .B2(new_n899_), .ZN(G69));
  XNOR2_X1  g728(.A(new_n666_), .B(KEYINPUT119), .ZN(new_n915_));
  NAND2_X1  g729(.A1(new_n815_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g730(.A1(new_n724_), .A2(new_n754_), .ZN(new_n917_));
  NAND3_X1  g731(.A1(new_n916_), .A2(new_n823_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n919_));
  NAND2_X1  g733(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND4_X1  g734(.A1(new_n916_), .A2(KEYINPUT120), .A3(new_n823_), .A4(new_n917_), .ZN(new_n921_));
  NAND2_X1  g735(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g736(.A1(new_n784_), .A2(new_n777_), .ZN(new_n923_));
  NOR3_X1   g737(.A1(new_n923_), .A2(new_n716_), .A3(new_n820_), .ZN(new_n924_));
  NAND3_X1  g738(.A1(new_n922_), .A2(new_n699_), .A3(new_n924_), .ZN(new_n925_));
  XOR2_X1   g739(.A(new_n343_), .B(KEYINPUT116), .Z(new_n926_));
  INV_X1    g740(.A(new_n926_), .ZN(new_n927_));
  NOR2_X1   g741(.A1(new_n556_), .A2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g742(.A1(new_n682_), .A2(G953), .ZN(new_n929_));
  OAI21_X1  g743(.A(new_n929_), .B1(new_n542_), .B2(new_n926_), .ZN(new_n930_));
  NOR2_X1   g744(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g745(.A(new_n931_), .ZN(new_n932_));
  NAND3_X1  g746(.A1(new_n925_), .A2(new_n281_), .A3(new_n932_), .ZN(new_n933_));
  NOR3_X1   g747(.A1(new_n687_), .A2(new_n691_), .A3(KEYINPUT79), .ZN(new_n934_));
  AOI21_X1  g748(.A(new_n697_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n935_));
  NOR2_X1   g749(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR3_X1   g750(.A1(new_n775_), .A2(new_n385_), .A3(new_n709_), .ZN(new_n937_));
  NAND3_X1  g751(.A1(new_n619_), .A2(new_n937_), .A3(new_n526_), .ZN(new_n938_));
  NAND3_X1  g752(.A1(new_n938_), .A2(new_n722_), .A3(new_n750_), .ZN(new_n939_));
  OAI21_X1  g753(.A(KEYINPUT117), .B1(new_n936_), .B2(new_n939_), .ZN(new_n940_));
  AND3_X1   g754(.A1(new_n938_), .A2(new_n722_), .A3(new_n750_), .ZN(new_n941_));
  INV_X1    g755(.A(KEYINPUT117), .ZN(new_n942_));
  NAND3_X1  g756(.A1(new_n941_), .A2(new_n699_), .A3(new_n942_), .ZN(new_n943_));
  AND3_X1   g757(.A1(new_n784_), .A2(new_n836_), .A3(new_n777_), .ZN(new_n944_));
  NAND3_X1  g758(.A1(new_n940_), .A2(new_n943_), .A3(new_n944_), .ZN(new_n945_));
  AOI211_X1 g759(.A(KEYINPUT118), .B(new_n932_), .C1(new_n945_), .C2(new_n277_), .ZN(new_n946_));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n947_));
  NAND2_X1  g761(.A1(new_n943_), .A2(new_n944_), .ZN(new_n948_));
  AOI21_X1  g762(.A(new_n942_), .B1(new_n941_), .B2(new_n699_), .ZN(new_n949_));
  OAI21_X1  g763(.A(new_n277_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g764(.A(new_n947_), .B1(new_n950_), .B2(new_n931_), .ZN(new_n951_));
  OAI21_X1  g765(.A(new_n933_), .B1(new_n946_), .B2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g766(.A(new_n281_), .B1(G227), .B2(G900), .ZN(new_n953_));
  INV_X1    g767(.A(new_n953_), .ZN(new_n954_));
  AND3_X1   g768(.A1(new_n952_), .A2(KEYINPUT121), .A3(new_n954_), .ZN(new_n955_));
  AOI21_X1  g769(.A(KEYINPUT121), .B1(new_n952_), .B2(new_n954_), .ZN(new_n956_));
  NOR2_X1   g770(.A1(new_n955_), .A2(new_n956_), .ZN(new_n957_));
  OAI211_X1 g771(.A(new_n953_), .B(new_n933_), .C1(new_n946_), .C2(new_n951_), .ZN(new_n958_));
  XNOR2_X1  g772(.A(new_n958_), .B(KEYINPUT122), .ZN(new_n959_));
  OAI21_X1  g773(.A(KEYINPUT123), .B1(new_n957_), .B2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g774(.A1(new_n952_), .A2(new_n954_), .ZN(new_n961_));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962_));
  NAND2_X1  g776(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g777(.A1(new_n952_), .A2(KEYINPUT121), .A3(new_n954_), .ZN(new_n964_));
  NAND2_X1  g778(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966_));
  XNOR2_X1  g780(.A(new_n958_), .B(new_n966_), .ZN(new_n967_));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n968_));
  NAND3_X1  g782(.A1(new_n965_), .A2(new_n967_), .A3(new_n968_), .ZN(new_n969_));
  NAND2_X1  g783(.A1(new_n960_), .A2(new_n969_), .ZN(G72));
  NAND2_X1  g784(.A1(new_n547_), .A2(new_n552_), .ZN(new_n971_));
  XNOR2_X1  g785(.A(new_n971_), .B(KEYINPUT124), .ZN(new_n972_));
  INV_X1    g786(.A(new_n972_), .ZN(new_n973_));
  NAND4_X1  g787(.A1(new_n844_), .A2(new_n922_), .A3(new_n699_), .A4(new_n924_), .ZN(new_n974_));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975_));
  AND3_X1   g789(.A1(new_n741_), .A2(new_n975_), .A3(new_n845_), .ZN(new_n976_));
  AOI21_X1  g790(.A(new_n975_), .B1(new_n741_), .B2(new_n845_), .ZN(new_n977_));
  NOR3_X1   g791(.A1(new_n974_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n978_));
  OAI21_X1  g792(.A(new_n973_), .B1(new_n978_), .B2(new_n573_), .ZN(new_n979_));
  NOR2_X1   g793(.A1(new_n973_), .A2(new_n573_), .ZN(new_n980_));
  INV_X1    g794(.A(new_n980_), .ZN(new_n981_));
  AOI21_X1  g795(.A(new_n981_), .B1(new_n850_), .B2(new_n843_), .ZN(new_n982_));
  OAI21_X1  g796(.A(new_n979_), .B1(new_n982_), .B2(KEYINPUT126), .ZN(new_n983_));
  AND2_X1   g797(.A1(new_n982_), .A2(KEYINPUT126), .ZN(new_n984_));
  OAI21_X1  g798(.A(new_n551_), .B1(new_n983_), .B2(new_n984_), .ZN(new_n985_));
  NAND2_X1  g799(.A1(new_n848_), .A2(new_n572_), .ZN(new_n986_));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987_));
  NAND3_X1  g801(.A1(new_n986_), .A2(new_n987_), .A3(new_n973_), .ZN(new_n988_));
  AOI21_X1  g802(.A(new_n573_), .B1(new_n850_), .B2(new_n843_), .ZN(new_n989_));
  OAI21_X1  g803(.A(KEYINPUT125), .B1(new_n989_), .B2(new_n972_), .ZN(new_n990_));
  OR2_X1    g804(.A1(new_n846_), .A2(new_n945_), .ZN(new_n991_));
  AOI21_X1  g805(.A(new_n551_), .B1(new_n991_), .B2(new_n980_), .ZN(new_n992_));
  NAND3_X1  g806(.A1(new_n988_), .A2(new_n990_), .A3(new_n992_), .ZN(new_n993_));
  AND3_X1   g807(.A1(new_n985_), .A2(new_n856_), .A3(new_n993_), .ZN(G57));
endmodule


